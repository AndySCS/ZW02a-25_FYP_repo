interface axi_rd_intf(
);

endinterface