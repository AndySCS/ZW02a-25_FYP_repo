class rf_output_transaction extends uvm_sequence_item;

    bit [31:0][31:0] rf_output;

    function new(string name = "rf_output_transaction");
       super.new(name);
    endfunction //new()

    `uvm_object_utils(rf_output_transaction)

endclass //top_tr extends superClass

