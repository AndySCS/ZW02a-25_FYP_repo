class mxu_output_monitor extends uvm_monitor;

    virtual mxu_intf mxu_if;
    uvm_analysis_port #(mxu_tr) ap;

    `uvm_component_utils(mxu_output_monitor)
    function new(string name = "mxu_output_monitor", uvm_component parent = null);
       super.new(name, parent);
    endfunction //new()
    
    extern virtual task build_phase(uvm_phase phase);
    extern virtual task main_phase(uvm_phase phase);
    
    extern virtual task collect_matrix_out(mxu_tr tr);

endclass //mxu_output_monitor extends superClass

task mxu_output_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual mxu_intf)::get(this, "", "mxu_if", mxu_if))begin
        `uvm_fatal("mxu_output_monitor", "mxu output_monitor fail to get mxu if")
    end
    ap = new("ap", this);
endtask

task mxu_output_monitor::main_phase(uvm_phase phase);
    mxu_tr tr;

    tr = new("tr");

    while (1) begin 
        this.collect_matrix_out(tr);
        ap.write(tr);
    end

endtask

task mxu_output_monitor::collect_matrix_out(mxu_tr tr);

    while(1)begin
        @(posedge mxu_if.clk);
        if(mxu_if.lsu_mxu_vld) break;
    end

    //tr.clear_result();
    @(posedge mxu_if.clk);
    wait(mxu_if.mxu_lsu_data_rdy) 
    tr.matrix_result[0][0] = $signed(mxu_if.mxu_lsu_int16_row0_data[15:0]);
    tr.matrix_result[0][1] = $signed(mxu_if.mxu_lsu_int16_row0_data[31:16]);
    tr.matrix_result[0][2] = $signed(mxu_if.mxu_lsu_int16_row0_data[47:32]);
    tr.matrix_result[0][3] = $signed(mxu_if.mxu_lsu_int16_row0_data[63:48]);
    tr.matrix_result[0][4] = $signed(mxu_if.mxu_lsu_int16_row0_data[79:64]);
    tr.matrix_result[0][5] = $signed(mxu_if.mxu_lsu_int16_row0_data[95:80]);
    tr.matrix_result[0][6] = $signed(mxu_if.mxu_lsu_int16_row0_data[111:96]);
    tr.matrix_result[0][7] = $signed(mxu_if.mxu_lsu_int16_row0_data[127:112]);
    tr.matrix_result[0][8] = $signed(mxu_if.mxu_lsu_int16_row0_data[143:128]);
    tr.matrix_result[0][9] = $signed(mxu_if.mxu_lsu_int16_row0_data[159:144]);
    tr.matrix_result[0][10] = $signed(mxu_if.mxu_lsu_int16_row0_data[175:160]);
    tr.matrix_result[0][11] = $signed(mxu_if.mxu_lsu_int16_row0_data[191:176]);
    tr.matrix_result[0][12] = $signed(mxu_if.mxu_lsu_int16_row0_data[207:192]);
    tr.matrix_result[0][13] = $signed(mxu_if.mxu_lsu_int16_row0_data[223:208]);
    tr.matrix_result[0][14] = $signed(mxu_if.mxu_lsu_int16_row0_data[239:224]);
    tr.matrix_result[0][15] = $signed(mxu_if.mxu_lsu_int16_row0_data[255:240]);
    tr.matrix_result[1][0] = $signed(mxu_if.mxu_lsu_int16_row1_data[15:0]);
    tr.matrix_result[1][1] = $signed(mxu_if.mxu_lsu_int16_row1_data[31:16]);
    tr.matrix_result[1][2] = $signed(mxu_if.mxu_lsu_int16_row1_data[47:32]);
    tr.matrix_result[1][3] = $signed(mxu_if.mxu_lsu_int16_row1_data[63:48]);
    tr.matrix_result[1][4] = $signed(mxu_if.mxu_lsu_int16_row1_data[79:64]);
    tr.matrix_result[1][5] = $signed(mxu_if.mxu_lsu_int16_row1_data[95:80]);
    tr.matrix_result[1][6] = $signed(mxu_if.mxu_lsu_int16_row1_data[111:96]);
    tr.matrix_result[1][7] = $signed(mxu_if.mxu_lsu_int16_row1_data[127:112]);
    tr.matrix_result[1][8] = $signed(mxu_if.mxu_lsu_int16_row1_data[143:128]);
    tr.matrix_result[1][9] = $signed(mxu_if.mxu_lsu_int16_row1_data[159:144]);
    tr.matrix_result[1][10] = $signed(mxu_if.mxu_lsu_int16_row1_data[175:160]);
    tr.matrix_result[1][11] = $signed(mxu_if.mxu_lsu_int16_row1_data[191:176]);
    tr.matrix_result[1][12] = $signed(mxu_if.mxu_lsu_int16_row1_data[207:192]);
    tr.matrix_result[1][13] = $signed(mxu_if.mxu_lsu_int16_row1_data[223:208]);
    tr.matrix_result[1][14] = $signed(mxu_if.mxu_lsu_int16_row1_data[239:224]);
    tr.matrix_result[1][15] = $signed(mxu_if.mxu_lsu_int16_row1_data[255:240]);
    tr.matrix_result[2][0] = $signed(mxu_if.mxu_lsu_int16_row2_data[15:0]);
    tr.matrix_result[2][1] = $signed(mxu_if.mxu_lsu_int16_row2_data[31:16]);
    tr.matrix_result[2][2] = $signed(mxu_if.mxu_lsu_int16_row2_data[47:32]);
    tr.matrix_result[2][3] = $signed(mxu_if.mxu_lsu_int16_row2_data[63:48]);
    tr.matrix_result[2][4] = $signed(mxu_if.mxu_lsu_int16_row2_data[79:64]);
    tr.matrix_result[2][5] = $signed(mxu_if.mxu_lsu_int16_row2_data[95:80]);
    tr.matrix_result[2][6] = $signed(mxu_if.mxu_lsu_int16_row2_data[111:96]);
    tr.matrix_result[2][7] = $signed(mxu_if.mxu_lsu_int16_row2_data[127:112]);
    tr.matrix_result[2][8] = $signed(mxu_if.mxu_lsu_int16_row2_data[143:128]);
    tr.matrix_result[2][9] = $signed(mxu_if.mxu_lsu_int16_row2_data[159:144]);
    tr.matrix_result[2][10] = $signed(mxu_if.mxu_lsu_int16_row2_data[175:160]);
    tr.matrix_result[2][11] = $signed(mxu_if.mxu_lsu_int16_row2_data[191:176]);
    tr.matrix_result[2][12] = $signed(mxu_if.mxu_lsu_int16_row2_data[207:192]);
    tr.matrix_result[2][13] = $signed(mxu_if.mxu_lsu_int16_row2_data[223:208]);
    tr.matrix_result[2][14] = $signed(mxu_if.mxu_lsu_int16_row2_data[239:224]);
    tr.matrix_result[2][15] = $signed(mxu_if.mxu_lsu_int16_row2_data[255:240]);
    tr.matrix_result[3][0] = $signed(mxu_if.mxu_lsu_int16_row3_data[15:0]);
    tr.matrix_result[3][1] = $signed(mxu_if.mxu_lsu_int16_row3_data[31:16]);
    tr.matrix_result[3][2] = $signed(mxu_if.mxu_lsu_int16_row3_data[47:32]);
    tr.matrix_result[3][3] = $signed(mxu_if.mxu_lsu_int16_row3_data[63:48]);
    tr.matrix_result[3][4] = $signed(mxu_if.mxu_lsu_int16_row3_data[79:64]);
    tr.matrix_result[3][5] = $signed(mxu_if.mxu_lsu_int16_row3_data[95:80]);
    tr.matrix_result[3][6] = $signed(mxu_if.mxu_lsu_int16_row3_data[111:96]);
    tr.matrix_result[3][7] = $signed(mxu_if.mxu_lsu_int16_row3_data[127:112]);
    tr.matrix_result[3][8] = $signed(mxu_if.mxu_lsu_int16_row3_data[143:128]);
    tr.matrix_result[3][9] = $signed(mxu_if.mxu_lsu_int16_row3_data[159:144]);
    tr.matrix_result[3][10] = $signed(mxu_if.mxu_lsu_int16_row3_data[175:160]);
    tr.matrix_result[3][11] = $signed(mxu_if.mxu_lsu_int16_row3_data[191:176]);
    tr.matrix_result[3][12] = $signed(mxu_if.mxu_lsu_int16_row3_data[207:192]);
    tr.matrix_result[3][13] = $signed(mxu_if.mxu_lsu_int16_row3_data[223:208]);
    tr.matrix_result[3][14] = $signed(mxu_if.mxu_lsu_int16_row3_data[239:224]);
    tr.matrix_result[3][15] = $signed(mxu_if.mxu_lsu_int16_row3_data[255:240]);
    tr.matrix_result[4][0] = $signed(mxu_if.mxu_lsu_int16_row4_data[15:0]);
    tr.matrix_result[4][1] = $signed(mxu_if.mxu_lsu_int16_row4_data[31:16]);
    tr.matrix_result[4][2] = $signed(mxu_if.mxu_lsu_int16_row4_data[47:32]);
    tr.matrix_result[4][3] = $signed(mxu_if.mxu_lsu_int16_row4_data[63:48]);
    tr.matrix_result[4][4] = $signed(mxu_if.mxu_lsu_int16_row4_data[79:64]);
    tr.matrix_result[4][5] = $signed(mxu_if.mxu_lsu_int16_row4_data[95:80]);
    tr.matrix_result[4][6] = $signed(mxu_if.mxu_lsu_int16_row4_data[111:96]);
    tr.matrix_result[4][7] = $signed(mxu_if.mxu_lsu_int16_row4_data[127:112]);
    tr.matrix_result[4][8] = $signed(mxu_if.mxu_lsu_int16_row4_data[143:128]);
    tr.matrix_result[4][9] = $signed(mxu_if.mxu_lsu_int16_row4_data[159:144]);
    tr.matrix_result[4][10] = $signed(mxu_if.mxu_lsu_int16_row4_data[175:160]);
    tr.matrix_result[4][11] = $signed(mxu_if.mxu_lsu_int16_row4_data[191:176]);
    tr.matrix_result[4][12] = $signed(mxu_if.mxu_lsu_int16_row4_data[207:192]);
    tr.matrix_result[4][13] = $signed(mxu_if.mxu_lsu_int16_row4_data[223:208]);
    tr.matrix_result[4][14] = $signed(mxu_if.mxu_lsu_int16_row4_data[239:224]);
    tr.matrix_result[4][15] = $signed(mxu_if.mxu_lsu_int16_row4_data[255:240]);
    tr.matrix_result[5][0] = $signed(mxu_if.mxu_lsu_int16_row5_data[15:0]);
    tr.matrix_result[5][1] = $signed(mxu_if.mxu_lsu_int16_row5_data[31:16]);
    tr.matrix_result[5][2] = $signed(mxu_if.mxu_lsu_int16_row5_data[47:32]);
    tr.matrix_result[5][3] = $signed(mxu_if.mxu_lsu_int16_row5_data[63:48]);
    tr.matrix_result[5][4] = $signed(mxu_if.mxu_lsu_int16_row5_data[79:64]);
    tr.matrix_result[5][5] = $signed(mxu_if.mxu_lsu_int16_row5_data[95:80]);
    tr.matrix_result[5][6] = $signed(mxu_if.mxu_lsu_int16_row5_data[111:96]);
    tr.matrix_result[5][7] = $signed(mxu_if.mxu_lsu_int16_row5_data[127:112]);
    tr.matrix_result[5][8] = $signed(mxu_if.mxu_lsu_int16_row5_data[143:128]);
    tr.matrix_result[5][9] = $signed(mxu_if.mxu_lsu_int16_row5_data[159:144]);
    tr.matrix_result[5][10] = $signed(mxu_if.mxu_lsu_int16_row5_data[175:160]);
    tr.matrix_result[5][11] = $signed(mxu_if.mxu_lsu_int16_row5_data[191:176]);
    tr.matrix_result[5][12] = $signed(mxu_if.mxu_lsu_int16_row5_data[207:192]);
    tr.matrix_result[5][13] = $signed(mxu_if.mxu_lsu_int16_row5_data[223:208]);
    tr.matrix_result[5][14] = $signed(mxu_if.mxu_lsu_int16_row5_data[239:224]);
    tr.matrix_result[5][15] = $signed(mxu_if.mxu_lsu_int16_row5_data[255:240]);
    tr.matrix_result[6][0] = $signed(mxu_if.mxu_lsu_int16_row6_data[15:0]);
    tr.matrix_result[6][1] = $signed(mxu_if.mxu_lsu_int16_row6_data[31:16]);
    tr.matrix_result[6][2] = $signed(mxu_if.mxu_lsu_int16_row6_data[47:32]);
    tr.matrix_result[6][3] = $signed(mxu_if.mxu_lsu_int16_row6_data[63:48]);
    tr.matrix_result[6][4] = $signed(mxu_if.mxu_lsu_int16_row6_data[79:64]);
    tr.matrix_result[6][5] = $signed(mxu_if.mxu_lsu_int16_row6_data[95:80]);
    tr.matrix_result[6][6] = $signed(mxu_if.mxu_lsu_int16_row6_data[111:96]);
    tr.matrix_result[6][7] = $signed(mxu_if.mxu_lsu_int16_row6_data[127:112]);
    tr.matrix_result[6][8] = $signed(mxu_if.mxu_lsu_int16_row6_data[143:128]);
    tr.matrix_result[6][9] = $signed(mxu_if.mxu_lsu_int16_row6_data[159:144]);
    tr.matrix_result[6][10] = $signed(mxu_if.mxu_lsu_int16_row6_data[175:160]);
    tr.matrix_result[6][11] = $signed(mxu_if.mxu_lsu_int16_row6_data[191:176]);
    tr.matrix_result[6][12] = $signed(mxu_if.mxu_lsu_int16_row6_data[207:192]);
    tr.matrix_result[6][13] = $signed(mxu_if.mxu_lsu_int16_row6_data[223:208]);
    tr.matrix_result[6][14] = $signed(mxu_if.mxu_lsu_int16_row6_data[239:224]);
    tr.matrix_result[6][15] = $signed(mxu_if.mxu_lsu_int16_row6_data[255:240]);
    tr.matrix_result[7][0] = $signed(mxu_if.mxu_lsu_int16_row7_data[15:0]);
    tr.matrix_result[7][1] = $signed(mxu_if.mxu_lsu_int16_row7_data[31:16]);
    tr.matrix_result[7][2] = $signed(mxu_if.mxu_lsu_int16_row7_data[47:32]);
    tr.matrix_result[7][3] = $signed(mxu_if.mxu_lsu_int16_row7_data[63:48]);
    tr.matrix_result[7][4] = $signed(mxu_if.mxu_lsu_int16_row7_data[79:64]);
    tr.matrix_result[7][5] = $signed(mxu_if.mxu_lsu_int16_row7_data[95:80]);
    tr.matrix_result[7][6] = $signed(mxu_if.mxu_lsu_int16_row7_data[111:96]);
    tr.matrix_result[7][7] = $signed(mxu_if.mxu_lsu_int16_row7_data[127:112]);
    tr.matrix_result[7][8] = $signed(mxu_if.mxu_lsu_int16_row7_data[143:128]);
    tr.matrix_result[7][9] = $signed(mxu_if.mxu_lsu_int16_row7_data[159:144]);
    tr.matrix_result[7][10] = $signed(mxu_if.mxu_lsu_int16_row7_data[175:160]);
    tr.matrix_result[7][11] = $signed(mxu_if.mxu_lsu_int16_row7_data[191:176]);
    tr.matrix_result[7][12] = $signed(mxu_if.mxu_lsu_int16_row7_data[207:192]);
    tr.matrix_result[7][13] = $signed(mxu_if.mxu_lsu_int16_row7_data[223:208]);
    tr.matrix_result[7][14] = $signed(mxu_if.mxu_lsu_int16_row7_data[239:224]);
    tr.matrix_result[7][15] = $signed(mxu_if.mxu_lsu_int16_row7_data[255:240]);
    tr.matrix_result[8][0] = $signed(mxu_if.mxu_lsu_int16_row8_data[15:0]);
    tr.matrix_result[8][1] = $signed(mxu_if.mxu_lsu_int16_row8_data[31:16]);
    tr.matrix_result[8][2] = $signed(mxu_if.mxu_lsu_int16_row8_data[47:32]);
    tr.matrix_result[8][3] = $signed(mxu_if.mxu_lsu_int16_row8_data[63:48]);
    tr.matrix_result[8][4] = $signed(mxu_if.mxu_lsu_int16_row8_data[79:64]);
    tr.matrix_result[8][5] = $signed(mxu_if.mxu_lsu_int16_row8_data[95:80]);
    tr.matrix_result[8][6] = $signed(mxu_if.mxu_lsu_int16_row8_data[111:96]);
    tr.matrix_result[8][7] = $signed(mxu_if.mxu_lsu_int16_row8_data[127:112]);
    tr.matrix_result[8][8] = $signed(mxu_if.mxu_lsu_int16_row8_data[143:128]);
    tr.matrix_result[8][9] = $signed(mxu_if.mxu_lsu_int16_row8_data[159:144]);
    tr.matrix_result[8][10] = $signed(mxu_if.mxu_lsu_int16_row8_data[175:160]);
    tr.matrix_result[8][11] = $signed(mxu_if.mxu_lsu_int16_row8_data[191:176]);
    tr.matrix_result[8][12] = $signed(mxu_if.mxu_lsu_int16_row8_data[207:192]);
    tr.matrix_result[8][13] = $signed(mxu_if.mxu_lsu_int16_row8_data[223:208]);
    tr.matrix_result[8][14] = $signed(mxu_if.mxu_lsu_int16_row8_data[239:224]);
    tr.matrix_result[8][15] = $signed(mxu_if.mxu_lsu_int16_row8_data[255:240]);
    tr.matrix_result[9][0] = $signed(mxu_if.mxu_lsu_int16_row9_data[15:0]);
    tr.matrix_result[9][1] = $signed(mxu_if.mxu_lsu_int16_row9_data[31:16]);
    tr.matrix_result[9][2] = $signed(mxu_if.mxu_lsu_int16_row9_data[47:32]);
    tr.matrix_result[9][3] = $signed(mxu_if.mxu_lsu_int16_row9_data[63:48]);
    tr.matrix_result[9][4] = $signed(mxu_if.mxu_lsu_int16_row9_data[79:64]);
    tr.matrix_result[9][5] = $signed(mxu_if.mxu_lsu_int16_row9_data[95:80]);
    tr.matrix_result[9][6] = $signed(mxu_if.mxu_lsu_int16_row9_data[111:96]);
    tr.matrix_result[9][7] = $signed(mxu_if.mxu_lsu_int16_row9_data[127:112]);
    tr.matrix_result[9][8] = $signed(mxu_if.mxu_lsu_int16_row9_data[143:128]);
    tr.matrix_result[9][9] = $signed(mxu_if.mxu_lsu_int16_row9_data[159:144]);
    tr.matrix_result[9][10] = $signed(mxu_if.mxu_lsu_int16_row9_data[175:160]);
    tr.matrix_result[9][11] = $signed(mxu_if.mxu_lsu_int16_row9_data[191:176]);
    tr.matrix_result[9][12] = $signed(mxu_if.mxu_lsu_int16_row9_data[207:192]);
    tr.matrix_result[9][13] = $signed(mxu_if.mxu_lsu_int16_row9_data[223:208]);
    tr.matrix_result[9][14] = $signed(mxu_if.mxu_lsu_int16_row9_data[239:224]);
    tr.matrix_result[9][15] = $signed(mxu_if.mxu_lsu_int16_row9_data[255:240]);
    tr.matrix_result[10][0] = $signed(mxu_if.mxu_lsu_int16_row10_data[15:0]);
    tr.matrix_result[10][1] = $signed(mxu_if.mxu_lsu_int16_row10_data[31:16]);
    tr.matrix_result[10][2] = $signed(mxu_if.mxu_lsu_int16_row10_data[47:32]);
    tr.matrix_result[10][3] = $signed(mxu_if.mxu_lsu_int16_row10_data[63:48]);
    tr.matrix_result[10][4] = $signed(mxu_if.mxu_lsu_int16_row10_data[79:64]);
    tr.matrix_result[10][5] = $signed(mxu_if.mxu_lsu_int16_row10_data[95:80]);
    tr.matrix_result[10][6] = $signed(mxu_if.mxu_lsu_int16_row10_data[111:96]);
    tr.matrix_result[10][7] = $signed(mxu_if.mxu_lsu_int16_row10_data[127:112]);
    tr.matrix_result[10][8] = $signed(mxu_if.mxu_lsu_int16_row10_data[143:128]);
    tr.matrix_result[10][9] = $signed(mxu_if.mxu_lsu_int16_row10_data[159:144]);
    tr.matrix_result[10][10] = $signed(mxu_if.mxu_lsu_int16_row10_data[175:160]);
    tr.matrix_result[10][11] = $signed(mxu_if.mxu_lsu_int16_row10_data[191:176]);
    tr.matrix_result[10][12] = $signed(mxu_if.mxu_lsu_int16_row10_data[207:192]);
    tr.matrix_result[10][13] = $signed(mxu_if.mxu_lsu_int16_row10_data[223:208]);
    tr.matrix_result[10][14] = $signed(mxu_if.mxu_lsu_int16_row10_data[239:224]);
    tr.matrix_result[10][15] = $signed(mxu_if.mxu_lsu_int16_row10_data[255:240]);
    tr.matrix_result[11][0] = $signed(mxu_if.mxu_lsu_int16_row11_data[15:0]);
    tr.matrix_result[11][1] = $signed(mxu_if.mxu_lsu_int16_row11_data[31:16]);
    tr.matrix_result[11][2] = $signed(mxu_if.mxu_lsu_int16_row11_data[47:32]);
    tr.matrix_result[11][3] = $signed(mxu_if.mxu_lsu_int16_row11_data[63:48]);
    tr.matrix_result[11][4] = $signed(mxu_if.mxu_lsu_int16_row11_data[79:64]);
    tr.matrix_result[11][5] = $signed(mxu_if.mxu_lsu_int16_row11_data[95:80]);
    tr.matrix_result[11][6] = $signed(mxu_if.mxu_lsu_int16_row11_data[111:96]);
    tr.matrix_result[11][7] = $signed(mxu_if.mxu_lsu_int16_row11_data[127:112]);
    tr.matrix_result[11][8] = $signed(mxu_if.mxu_lsu_int16_row11_data[143:128]);
    tr.matrix_result[11][9] = $signed(mxu_if.mxu_lsu_int16_row11_data[159:144]);
    tr.matrix_result[11][10] = $signed(mxu_if.mxu_lsu_int16_row11_data[175:160]);
    tr.matrix_result[11][11] = $signed(mxu_if.mxu_lsu_int16_row11_data[191:176]);
    tr.matrix_result[11][12] = $signed(mxu_if.mxu_lsu_int16_row11_data[207:192]);
    tr.matrix_result[11][13] = $signed(mxu_if.mxu_lsu_int16_row11_data[223:208]);
    tr.matrix_result[11][14] = $signed(mxu_if.mxu_lsu_int16_row11_data[239:224]);
    tr.matrix_result[11][15] = $signed(mxu_if.mxu_lsu_int16_row11_data[255:240]);
    tr.matrix_result[12][0] = $signed(mxu_if.mxu_lsu_int16_row12_data[15:0]);
    tr.matrix_result[12][1] = $signed(mxu_if.mxu_lsu_int16_row12_data[31:16]);
    tr.matrix_result[12][2] = $signed(mxu_if.mxu_lsu_int16_row12_data[47:32]);
    tr.matrix_result[12][3] = $signed(mxu_if.mxu_lsu_int16_row12_data[63:48]);
    tr.matrix_result[12][4] = $signed(mxu_if.mxu_lsu_int16_row12_data[79:64]);
    tr.matrix_result[12][5] = $signed(mxu_if.mxu_lsu_int16_row12_data[95:80]);
    tr.matrix_result[12][6] = $signed(mxu_if.mxu_lsu_int16_row12_data[111:96]);
    tr.matrix_result[12][7] = $signed(mxu_if.mxu_lsu_int16_row12_data[127:112]);
    tr.matrix_result[12][8] = $signed(mxu_if.mxu_lsu_int16_row12_data[143:128]);
    tr.matrix_result[12][9] = $signed(mxu_if.mxu_lsu_int16_row12_data[159:144]);
    tr.matrix_result[12][10] = $signed(mxu_if.mxu_lsu_int16_row12_data[175:160]);
    tr.matrix_result[12][11] = $signed(mxu_if.mxu_lsu_int16_row12_data[191:176]);
    tr.matrix_result[12][12] = $signed(mxu_if.mxu_lsu_int16_row12_data[207:192]);
    tr.matrix_result[12][13] = $signed(mxu_if.mxu_lsu_int16_row12_data[223:208]);
    tr.matrix_result[12][14] = $signed(mxu_if.mxu_lsu_int16_row12_data[239:224]);
    tr.matrix_result[12][15] = $signed(mxu_if.mxu_lsu_int16_row12_data[255:240]);
    tr.matrix_result[13][0] = $signed(mxu_if.mxu_lsu_int16_row13_data[15:0]);
    tr.matrix_result[13][1] = $signed(mxu_if.mxu_lsu_int16_row13_data[31:16]);
    tr.matrix_result[13][2] = $signed(mxu_if.mxu_lsu_int16_row13_data[47:32]);
    tr.matrix_result[13][3] = $signed(mxu_if.mxu_lsu_int16_row13_data[63:48]);
    tr.matrix_result[13][4] = $signed(mxu_if.mxu_lsu_int16_row13_data[79:64]);
    tr.matrix_result[13][5] = $signed(mxu_if.mxu_lsu_int16_row13_data[95:80]);
    tr.matrix_result[13][6] = $signed(mxu_if.mxu_lsu_int16_row13_data[111:96]);
    tr.matrix_result[13][7] = $signed(mxu_if.mxu_lsu_int16_row13_data[127:112]);
    tr.matrix_result[13][8] = $signed(mxu_if.mxu_lsu_int16_row13_data[143:128]);
    tr.matrix_result[13][9] = $signed(mxu_if.mxu_lsu_int16_row13_data[159:144]);
    tr.matrix_result[13][10] = $signed(mxu_if.mxu_lsu_int16_row13_data[175:160]);
    tr.matrix_result[13][11] = $signed(mxu_if.mxu_lsu_int16_row13_data[191:176]);
    tr.matrix_result[13][12] = $signed(mxu_if.mxu_lsu_int16_row13_data[207:192]);
    tr.matrix_result[13][13] = $signed(mxu_if.mxu_lsu_int16_row13_data[223:208]);
    tr.matrix_result[13][14] = $signed(mxu_if.mxu_lsu_int16_row13_data[239:224]);
    tr.matrix_result[13][15] = $signed(mxu_if.mxu_lsu_int16_row13_data[255:240]);
    tr.matrix_result[14][0] = $signed(mxu_if.mxu_lsu_int16_row14_data[15:0]);
    tr.matrix_result[14][1] = $signed(mxu_if.mxu_lsu_int16_row14_data[31:16]);
    tr.matrix_result[14][2] = $signed(mxu_if.mxu_lsu_int16_row14_data[47:32]);
    tr.matrix_result[14][3] = $signed(mxu_if.mxu_lsu_int16_row14_data[63:48]);
    tr.matrix_result[14][4] = $signed(mxu_if.mxu_lsu_int16_row14_data[79:64]);
    tr.matrix_result[14][5] = $signed(mxu_if.mxu_lsu_int16_row14_data[95:80]);
    tr.matrix_result[14][6] = $signed(mxu_if.mxu_lsu_int16_row14_data[111:96]);
    tr.matrix_result[14][7] = $signed(mxu_if.mxu_lsu_int16_row14_data[127:112]);
    tr.matrix_result[14][8] = $signed(mxu_if.mxu_lsu_int16_row14_data[143:128]);
    tr.matrix_result[14][9] = $signed(mxu_if.mxu_lsu_int16_row14_data[159:144]);
    tr.matrix_result[14][10] = $signed(mxu_if.mxu_lsu_int16_row14_data[175:160]);
    tr.matrix_result[14][11] = $signed(mxu_if.mxu_lsu_int16_row14_data[191:176]);
    tr.matrix_result[14][12] = $signed(mxu_if.mxu_lsu_int16_row14_data[207:192]);
    tr.matrix_result[14][13] = $signed(mxu_if.mxu_lsu_int16_row14_data[223:208]);
    tr.matrix_result[14][14] = $signed(mxu_if.mxu_lsu_int16_row14_data[239:224]);
    tr.matrix_result[14][15] = $signed(mxu_if.mxu_lsu_int16_row14_data[255:240]);
    tr.matrix_result[15][0] = $signed(mxu_if.mxu_lsu_int16_row15_data[15:0]);
    tr.matrix_result[15][1] = $signed(mxu_if.mxu_lsu_int16_row15_data[31:16]);
    tr.matrix_result[15][2] = $signed(mxu_if.mxu_lsu_int16_row15_data[47:32]);
    tr.matrix_result[15][3] = $signed(mxu_if.mxu_lsu_int16_row15_data[63:48]);
    tr.matrix_result[15][4] = $signed(mxu_if.mxu_lsu_int16_row15_data[79:64]);
    tr.matrix_result[15][5] = $signed(mxu_if.mxu_lsu_int16_row15_data[95:80]);
    tr.matrix_result[15][6] = $signed(mxu_if.mxu_lsu_int16_row15_data[111:96]);
    tr.matrix_result[15][7] = $signed(mxu_if.mxu_lsu_int16_row15_data[127:112]);
    tr.matrix_result[15][8] = $signed(mxu_if.mxu_lsu_int16_row15_data[143:128]);
    tr.matrix_result[15][9] = $signed(mxu_if.mxu_lsu_int16_row15_data[159:144]);
    tr.matrix_result[15][10] = $signed(mxu_if.mxu_lsu_int16_row15_data[175:160]);
    tr.matrix_result[15][11] = $signed(mxu_if.mxu_lsu_int16_row15_data[191:176]);
    tr.matrix_result[15][12] = $signed(mxu_if.mxu_lsu_int16_row15_data[207:192]);
    tr.matrix_result[15][13] = $signed(mxu_if.mxu_lsu_int16_row15_data[223:208]);
    tr.matrix_result[15][14] = $signed(mxu_if.mxu_lsu_int16_row15_data[239:224]);
    tr.matrix_result[15][15] = $signed(mxu_if.mxu_lsu_int16_row15_data[255:240]);

endtask
