interface start_if;
    
endinterface