class tc_base extends uvm_test;

    env tc_env;

    function new(string name = "tc_base", uvm_component parent = null);
        super.new(name, parent);
    endfunction //new()

    extern function void build_phase(uvm_phase phase);
    extern function void connect_phase(uvm_phase phase);
    extern task reset_phase(uvm_phase phase);
    extern function void report_phase(uvm_phase phase);

    `uvm_component_utils(tc_base)

endclass

function void tc_base::build_phase(uvm_phase phase);
    `uvm_info(get_name(), "build phase begins", UVM_LOW);
    super.build_phase(phase);
    tc_env = env::type_id::create("tc_env", this);
    `uvm_info(get_name(), "build phase ends", UVM_LOW);
endfunction

function void tc_base::connect_phase(uvm_phase phase);
    `uvm_info(get_name(), "connect phase begins", UVM_LOW);
    super.connect_phase(phase);
    `uvm_info(get_name(), "connect phase ends", UVM_LOW);
endfunction

task tc_base::reset_phase(uvm_phase phase);
    `uvm_info(get_name(), "reset phase begins", UVM_LOW);
    super.reset_phase(phase);
    `uvm_info(get_name(), "reset phase ends", UVM_LOW);
endtask

function void tc_base::report_phase(uvm_phase phase);

    int err_num;    

    uvm_report_server server;
    super.report_phase(phase);

    server = get_report_server();
    err_num = server.get_severity_count(UVM_ERROR);

    if(err_num > 0) $display("TC ERROR");
    else $display("TC PASS");

endfunction
