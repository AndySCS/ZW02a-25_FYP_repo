module sixteen_ff(
    in,
    out
);

    input [15:0] in;
    output [15:0] out;

    assign out = in[0] ?  16'b0000_0000_0000_0001
               : in[1] ?  16'b0000_0000_0000_0010
               : in[2] ?  16'b0000_0000_0000_0100
               : in[3] ?  16'b0000_0000_0000_1000
               : in[4] ?  16'b0000_0000_0001_0000
               : in[5] ?  16'b0000_0000_0010_0000
               : in[6] ?  16'b0000_0000_0100_0000
               : in[7] ?  16'b0000_0000_1000_0000
               : in[8] ?  16'b0000_0001_0000_0000
               : in[9] ?  16'b0000_0010_0000_0000
               : in[10] ? 16'b0000_0100_0000_0000
               : in[11] ? 16'b0000_1000_0000_0000
               : in[12] ? 16'b0001_0000_0000_0000
               : in[13] ? 16'b0010_0000_0000_0000
               : in[14] ? 16'b0100_0000_0000_0000
               : in[15] ? 16'b1000_0000_0000_0000
               : 16'h0000;

endmodule