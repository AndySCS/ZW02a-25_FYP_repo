module dec5to32(
    in,
    out
);
    input [4:0] in;
    output reg [31:0] out;

    always @(*) begin
        case (in)
            5'd0 : out <= 16'b0000_0000_0000_0000_0000_0000_0000_0001;
            5'd1 : out <= 16'b0000_0000_0000_0000_0000_0000_0000_0010;
            5'd2 : out <= 16'b0000_0000_0000_0000_0000_0000_0000_0100;
            5'd3 : out <= 16'b0000_0000_0000_0000_0000_0000_0000_1000;
            5'd4 : out <= 16'b0000_0000_0000_0000_0000_0000_0001_0000;
            5'd5 : out <= 16'b0000_0000_0000_0000_0000_0000_0010_0000;
            5'd6 : out <= 16'b0000_0000_0000_0000_0000_0000_0100_0000;
            5'd7 : out <= 16'b0000_0000_0000_0000_0000_0000_1000_0000;
            5'd8 : out <= 16'b0000_0000_0000_0000_0000_0001_0000_0000;
            5'd9 : out <= 16'b0000_0000_0000_0000_0000_0010_0000_0000;
            5'd10: out <= 16'b0000_0000_0000_0000_0000_0100_0000_0000;
            5'd11: out <= 16'b0000_0000_0000_0000_0000_1000_0000_0000;
            5'd12: out <= 16'b0000_0000_0000_0000_0001_0000_0000_0000;
            5'd13: out <= 16'b0000_0000_0000_0000_0010_0000_0000_0000;
            5'd14: out <= 16'b0000_0000_0000_0000_0100_0000_0000_0000;
            5'd15: out <= 16'b0000_0000_0000_0000_1000_0000_0000_0000;
            5'd16: out <= 16'b0000_0000_0000_0001_0000_0000_0000_0000;
            5'd17: out <= 16'b0000_0000_0000_0010_0000_0000_0000_0000;
            5'd18: out <= 16'b0000_0000_0000_0100_0000_0000_0000_0000;
            5'd19: out <= 16'b0000_0000_0000_1000_0000_0000_0000_0000;
            5'd20: out <= 16'b0000_0000_0001_0000_0000_0000_0000_0000;
            5'd21: out <= 16'b0000_0000_0010_0000_0000_0000_0000_0000;
            5'd22: out <= 16'b0000_0000_0100_0000_0000_0000_0000_0000;
            5'd23: out <= 16'b0000_0000_1000_0000_0000_0000_0000_0000;
            5'd24: out <= 16'b0000_0001_0000_0000_0000_0000_0000_0000;
            5'd25: out <= 16'b0000_0010_0000_0000_0000_0000_0000_0000;
            5'd26: out <= 16'b0000_0100_0000_0000_0000_0000_0000_0000;
            5'd27: out <= 16'b0000_1000_0000_0000_0000_0000_0000_0000;
            5'd28: out <= 16'b0001_0000_0000_0000_0000_0000_0000_0000;
            5'd29: out <= 16'b0010_0000_0000_0000_0000_0000_0000_0000;
            5'd30: out <= 16'b0100_0000_0000_0000_0000_0000_0000_0000;
            5'd31: out <= 16'b1000_0000_0000_0000_0000_0000_0000_0000;
            default: out <= 32'hxxxx_xxxx;
        endcase
    end

endmodule