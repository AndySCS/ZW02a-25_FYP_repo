module mxu (
    clk,
    rst_n,
    lsu_mxu_vld,
    lsu_mxu_clr,
    lsu_mxu_iram_vld,
    lsu_mxu_iram_pld,
    lsu_mxu_wram_vld,
    lsu_mxu_wram_pld,
    lsu_mxu_pool_vld,
    lsu_mxu_pool_size,
    lsu_mxu_act_vld,
    lsu_mxu_act_type,
    lsu_mxu_wfi,
    mxu_lsu_int8_row0_data,
    mxu_lsu_int16_row0_data,
    mxu_lsu_int8_row1_data,
    mxu_lsu_int16_row1_data,
    mxu_lsu_int8_row2_data,
    mxu_lsu_int16_row2_data,
    mxu_lsu_int8_row3_data,
    mxu_lsu_int16_row3_data,
    mxu_lsu_int8_row4_data,
    mxu_lsu_int16_row4_data,
    mxu_lsu_int8_row5_data,
    mxu_lsu_int16_row5_data,
    mxu_lsu_int8_row6_data,
    mxu_lsu_int16_row6_data,
    mxu_lsu_int8_row7_data,
    mxu_lsu_int16_row7_data,
    mxu_lsu_int8_row8_data,
    mxu_lsu_int16_row8_data,
    mxu_lsu_int8_row9_data,
    mxu_lsu_int16_row9_data,
    mxu_lsu_int8_row10_data,
    mxu_lsu_int16_row10_data,
    mxu_lsu_int8_row11_data,
    mxu_lsu_int16_row11_data,
    mxu_lsu_int8_row12_data,
    mxu_lsu_int16_row12_data,
    mxu_lsu_int8_row13_data,
    mxu_lsu_int16_row13_data,
    mxu_lsu_int8_row14_data,
    mxu_lsu_int16_row14_data,
    mxu_lsu_int8_row15_data,
    mxu_lsu_int16_row15_data,
    mxu_lsu_data_rdy,
    mxu_lsu_rdy
);
   
    input clk;
    input rst_n;
    input lsu_mxu_vld;
    input lsu_mxu_clr;
    input [15:0] lsu_mxu_iram_vld;
    input [127:0] lsu_mxu_iram_pld;
    input [15:0] lsu_mxu_wram_vld;
    input [127:0] lsu_mxu_wram_pld;
    input lsu_mxu_pool_vld;
    input [1:0] lsu_mxu_pool_size;
    input lsu_mxu_act_vld;
    input [1:0] lsu_mxu_act_type;
    input lsu_mxu_wfi;
    output [127:0] mxu_lsu_int8_row0_data;
    output [255:0] mxu_lsu_int16_row0_data;
    output [127:0] mxu_lsu_int8_row1_data;
    output [255:0] mxu_lsu_int16_row1_data;
    output [127:0] mxu_lsu_int8_row2_data;
    output [255:0] mxu_lsu_int16_row2_data;
    output [127:0] mxu_lsu_int8_row3_data;
    output [255:0] mxu_lsu_int16_row3_data;
    output [127:0] mxu_lsu_int8_row4_data;
    output [255:0] mxu_lsu_int16_row4_data;
    output [127:0] mxu_lsu_int8_row5_data;
    output [255:0] mxu_lsu_int16_row5_data;
    output [127:0] mxu_lsu_int8_row6_data;
    output [255:0] mxu_lsu_int16_row6_data;
    output [127:0] mxu_lsu_int8_row7_data;
    output [255:0] mxu_lsu_int16_row7_data;
    output [127:0] mxu_lsu_int8_row8_data;
    output [255:0] mxu_lsu_int16_row8_data;
    output [127:0] mxu_lsu_int8_row9_data;
    output [255:0] mxu_lsu_int16_row9_data;
    output [127:0] mxu_lsu_int8_row10_data;
    output [255:0] mxu_lsu_int16_row10_data;
    output [127:0] mxu_lsu_int8_row11_data;
    output [255:0] mxu_lsu_int16_row11_data;
    output [127:0] mxu_lsu_int8_row12_data;
    output [255:0] mxu_lsu_int16_row12_data;
    output [127:0] mxu_lsu_int8_row13_data;
    output [255:0] mxu_lsu_int16_row13_data;
    output [127:0] mxu_lsu_int8_row14_data;
    output [255:0] mxu_lsu_int16_row14_data;
    output [127:0] mxu_lsu_int8_row15_data;
    output [255:0] mxu_lsu_int16_row15_data;
    output mxu_lsu_data_rdy;
    output mxu_lsu_rdy;

    wire lsu_mxu_vld_qual;
    wire mxu_vld;
    wire mxu_vld_nxt;
    wire mxu_done;

    wire acc_clr;

    wire [15:0] c1_vld [15:0];
    wire [127:0] c1_data [15:0];

    wire mxu_act_vld;
    wire [15:0] act_vld [15:0];
    wire [255:0] act_data [15:0];
    wire act_busy;

    wire mxu_conv_awake_cnt_en;
    wire [2:0] mxu_conv_awake_cnt;   
    wire [2:0] mxu_conv_awake_cnt_nxt;
    wire [2:0] mxu_conv_awake_cnt_minus;

    
    wire [15:0] sys_arr_row0_load_vld;
    wire [127:0] sys_arr_row0_load_data;

    wire [15:0] sys_arr_row1_load_vld;
    wire [127:0] sys_arr_row1_load_data;

    wire [15:0] sys_arr_row2_load_vld;
    wire [127:0] sys_arr_row2_load_data;

    wire [15:0] sys_arr_row3_load_vld;
    wire [127:0] sys_arr_row3_load_data;

    wire [15:0] sys_arr_row4_load_vld;
    wire [127:0] sys_arr_row4_load_data;

    wire [15:0] sys_arr_row5_load_vld;
    wire [127:0] sys_arr_row5_load_data;

    wire [15:0] sys_arr_row6_load_vld;
    wire [127:0] sys_arr_row6_load_data;

    wire [15:0] sys_arr_row7_load_vld;
    wire [127:0] sys_arr_row7_load_data;

    wire [15:0] sys_arr_row8_load_vld;
    wire [127:0] sys_arr_row8_load_data;

    wire [15:0] sys_arr_row9_load_vld;
    wire [127:0] sys_arr_row9_load_data;

    wire [15:0] sys_arr_row10_load_vld;
    wire [127:0] sys_arr_row10_load_data;

    wire [15:0] sys_arr_row11_load_vld;
    wire [127:0] sys_arr_row11_load_data;

    wire [15:0] sys_arr_row12_load_vld;
    wire [127:0] sys_arr_row12_load_data;

    wire [15:0] sys_arr_row13_load_vld;
    wire [127:0] sys_arr_row13_load_data;

    wire [15:0] sys_arr_row14_load_vld;
    wire [127:0] sys_arr_row14_load_data;

    wire [15:0] sys_arr_row15_load_vld;
    wire [127:0] sys_arr_row15_load_data;

    wire [15:0] sys_arr_row16_load_vld;
    wire [127:0] sys_arr_row16_load_data;

    wire [15:0] sys_arr_row_data_rdy;

    assign sys_arr_row0_load_vld = act_vld[0];
    assign sys_arr_row0_load_data = act_data[0];
    assign sys_arr_row_data_rdy[0] = ~(|c1_vld[0]) & ~(|sys_arr_row0_load_vld) & ~(|pe_doing[0]);
    assign sys_arr_row1_load_vld = act_vld[1];
    assign sys_arr_row1_load_data = act_data[1];
    assign sys_arr_row_data_rdy[1] = ~(|c1_vld[1]) & ~(|sys_arr_row1_load_vld) & ~(|pe_doing[1]);
    assign sys_arr_row2_load_vld = act_vld[2];
    assign sys_arr_row2_load_data = act_data[2];
    assign sys_arr_row_data_rdy[2] = ~(|c1_vld[2]) & ~(|sys_arr_row2_load_vld) & ~(|pe_doing[2]);
    assign sys_arr_row3_load_vld = act_vld[3];
    assign sys_arr_row3_load_data = act_data[3];
    assign sys_arr_row_data_rdy[3] = ~(|c1_vld[3]) & ~(|sys_arr_row3_load_vld) & ~(|pe_doing[3]);
    assign sys_arr_row4_load_vld = act_vld[4];
    assign sys_arr_row4_load_data = act_data[4];
    assign sys_arr_row_data_rdy[4] = ~(|c1_vld[4]) & ~(|sys_arr_row4_load_vld) & ~(|pe_doing[4]);
    assign sys_arr_row5_load_vld = act_vld[5];
    assign sys_arr_row5_load_data = act_data[5];
    assign sys_arr_row_data_rdy[5] = ~(|c1_vld[5]) & ~(|sys_arr_row5_load_vld) & ~(|pe_doing[5]);
    assign sys_arr_row6_load_vld = act_vld[6];
    assign sys_arr_row6_load_data = act_data[6];
    assign sys_arr_row_data_rdy[6] = ~(|c1_vld[6]) & ~(|sys_arr_row6_load_vld) & ~(|pe_doing[6]);
    assign sys_arr_row7_load_vld = act_vld[7];
    assign sys_arr_row7_load_data = act_data[7];
    assign sys_arr_row_data_rdy[7] = ~(|c1_vld[7]) & ~(|sys_arr_row7_load_vld) & ~(|pe_doing[7]);
    assign sys_arr_row8_load_vld = act_vld[8];
    assign sys_arr_row8_load_data = act_data[8];
    assign sys_arr_row_data_rdy[8] = ~(|c1_vld[8]) & ~(|sys_arr_row8_load_vld) & ~(|pe_doing[8]);
    assign sys_arr_row9_load_vld = act_vld[9];
    assign sys_arr_row9_load_data = act_data[9];
    assign sys_arr_row_data_rdy[9] = ~(|c1_vld[9]) & ~(|sys_arr_row9_load_vld) & ~(|pe_doing[9]);
    assign sys_arr_row10_load_vld = act_vld[10];
    assign sys_arr_row10_load_data = act_data[10];
    assign sys_arr_row_data_rdy[10] = ~(|c1_vld[10]) & ~(|sys_arr_row10_load_vld) & ~(|pe_doing[10]);
    assign sys_arr_row11_load_vld = act_vld[11];
    assign sys_arr_row11_load_data = act_data[11];
    assign sys_arr_row_data_rdy[11] = ~(|c1_vld[11]) & ~(|sys_arr_row11_load_vld) & ~(|pe_doing[11]);
    assign sys_arr_row12_load_vld = act_vld[12];
    assign sys_arr_row12_load_data = act_data[12];
    assign sys_arr_row_data_rdy[12] = ~(|c1_vld[12]) & ~(|sys_arr_row12_load_vld) & ~(|pe_doing[12]);
    assign sys_arr_row13_load_vld = act_vld[13];
    assign sys_arr_row13_load_data = act_data[13];
    assign sys_arr_row_data_rdy[13] = ~(|c1_vld[13]) & ~(|sys_arr_row13_load_vld) & ~(|pe_doing[13]);
    assign sys_arr_row14_load_vld = act_vld[14];
    assign sys_arr_row14_load_data = act_data[14];
    assign sys_arr_row_data_rdy[14] = ~(|c1_vld[14]) & ~(|sys_arr_row14_load_vld) & ~(|pe_doing[14]);
    assign sys_arr_row15_load_vld = act_vld[15];
    assign sys_arr_row15_load_data = act_data[15];
    assign sys_arr_row_data_rdy[15] = ~(|c1_vld[15]) & ~(|sys_arr_row15_load_vld) & ~(|pe_doing[15]);
    assign sys_arr_row16_load_vld = act_vld[16];
    assign sys_arr_row16_load_data = act_data[16];
    assign sys_arr_row_data_rdy[16] = ~(|c1_vld[16]) & ~(|sys_arr_row16_load_vld) & ~(|pe_doing[16]);

    assign lsu_mxu_vld_qual = lsu_mxu_vld & mxu_lsu_rdy;
    assign mxu_vld_nxt = lsu_mxu_vld_qual | mxu_vld & ~mxu_done;

    assign mxu_done =  ~(|mxu_conv_awake_cnt_minus) & (|sys_arr_row_data_rdy);
    assign mxu_lsu_rdy = mxu_done | ~mxu_vld;

    assign mxu_lsu_data_rdy =  (|sys_arr_row_data_rdy) & ~act_busy ;

    DFFR #(.WIDTH(1))
    ff_mxu_vld(
        .clk(clk),
        .rst_n(rst_n),
        .d(mxu_vld_nxt),
        .q(mxu_vld)
    );

    assign acc_clr_qual = lsu_mxu_clr & lsu_mxu_vld_qual;
    assign mxu_act_vld = lsu_mxu_act_vld & lsu_mxu_vld_qual;

    assign mxu_conv_awake_cnt_en = (|mxu_conv_awake_cnt) | lsu_mxu_vld_qual;
    assign mxu_conv_awake_cnt_minus = mxu_conv_awake_cnt - 3'b1;
    assign mxu_conv_awake_cnt_nxt = lsu_mxu_clr ? 3'b111 : mxu_conv_awake_cnt_minus;

    DFFRE #(.WIDTH(3))
    ff_mxu_conv_awake_cnt(
        .clk(clk),
        .rst_n(rst_n),
        .en(mxu_conv_awake_cnt_en),
        .d(mxu_conv_awake_cnt_nxt),
        .q(mxu_conv_awake_cnt)
    );



    wire [15:0] sys_arr_row0_vld;
    wire [127:0] sys_arr_row0_data;
    wire [15:0] sys_arr_row1_vld;
    wire [127:0] sys_arr_row1_data;
    wire [15:0] sys_arr_row2_vld;
    wire [127:0] sys_arr_row2_data;
    wire [15:0] sys_arr_row3_vld;
    wire [127:0] sys_arr_row3_data;
    wire [15:0] sys_arr_row4_vld;
    wire [127:0] sys_arr_row4_data;
    wire [15:0] sys_arr_row5_vld;
    wire [127:0] sys_arr_row5_data;
    wire [15:0] sys_arr_row6_vld;
    wire [127:0] sys_arr_row6_data;
    wire [15:0] sys_arr_row7_vld;
    wire [127:0] sys_arr_row7_data;
    wire [15:0] sys_arr_row8_vld;
    wire [127:0] sys_arr_row8_data;
    wire [15:0] sys_arr_row9_vld;
    wire [127:0] sys_arr_row9_data;
    wire [15:0] sys_arr_row10_vld;
    wire [127:0] sys_arr_row10_data;
    wire [15:0] sys_arr_row11_vld;
    wire [127:0] sys_arr_row11_data;
    wire [15:0] sys_arr_row12_vld;
    wire [127:0] sys_arr_row12_data;
    wire [15:0] sys_arr_row13_vld;
    wire [127:0] sys_arr_row13_data;
    wire [15:0] sys_arr_row14_vld;
    wire [127:0] sys_arr_row14_data;
    wire [15:0] sys_arr_row15_vld;
    wire [127:0] sys_arr_row15_data;
    wire [15:0] sys_arr_row16_vld;
    wire [127:0] sys_arr_row16_data;

    wire [15:0] sys_arr_col0_vld;
    wire [127:0] sys_arr_col0_data;
    wire [15:0] sys_arr_col1_vld;
    wire [127:0] sys_arr_col1_data;
    wire [15:0] sys_arr_col2_vld;
    wire [127:0] sys_arr_col2_data;
    wire [15:0] sys_arr_col3_vld;
    wire [127:0] sys_arr_col3_data;
    wire [15:0] sys_arr_col4_vld;
    wire [127:0] sys_arr_col4_data;
    wire [15:0] sys_arr_col5_vld;
    wire [127:0] sys_arr_col5_data;
    wire [15:0] sys_arr_col6_vld;
    wire [127:0] sys_arr_col6_data;
    wire [15:0] sys_arr_col7_vld;
    wire [127:0] sys_arr_col7_data;
    wire [15:0] sys_arr_col8_vld;
    wire [127:0] sys_arr_col8_data;
    wire [15:0] sys_arr_col9_vld;
    wire [127:0] sys_arr_col9_data;
    wire [15:0] sys_arr_col10_vld;
    wire [127:0] sys_arr_col10_data;
    wire [15:0] sys_arr_col11_vld;
    wire [127:0] sys_arr_col11_data;
    wire [15:0] sys_arr_col12_vld;
    wire [127:0] sys_arr_col12_data;
    wire [15:0] sys_arr_col13_vld;
    wire [127:0] sys_arr_col13_data;
    wire [15:0] sys_arr_col14_vld;
    wire [127:0] sys_arr_col14_data;
    wire [15:0] sys_arr_col15_vld;
    wire [127:0] sys_arr_col15_data;
    wire [15:0] sys_arr_col16_vld;
    wire [127:0] sys_arr_col16_data;

    wire [15:0] pe_doing [15:0];

    assign sys_arr_row0_vld  = lsu_mxu_iram_vld;
    assign sys_arr_row0_data = lsu_mxu_iram_pld;
    assign sys_arr_col0_vld  = lsu_mxu_wram_vld;
    assign sys_arr_col0_data = lsu_mxu_wram_pld;

    pe u_pe_row0_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[0]),
        .in0_data(sys_arr_row0_data[7:0]),
        .in1_vld(sys_arr_col0_vld[0]),
        .in1_data(sys_arr_col0_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[0]),
        .out0_data(sys_arr_row1_data[7:0]),
        .out1_vld(sys_arr_col1_vld[0]),
        .out1_data(sys_arr_col1_data[7:0]),
        .pe_doing(pe_doing[0][0]),
        .c1_vld(c1_vld[0][0]),
        .c1_data(c1_data[0][7:0])
    );
    
    pe u_pe_row0_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[1]),
        .in0_data(sys_arr_row0_data[15:8]),
        .in1_vld(sys_arr_col1_vld[0]),
        .in1_data(sys_arr_col1_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[1]),
        .out0_data(sys_arr_row1_data[15:8]),
        .out1_vld(sys_arr_col2_vld[0]),
        .out1_data(sys_arr_col2_data[7:0]),
        .pe_doing(pe_doing[0][1]),
        .c1_vld(c1_vld[0][1]),
        .c1_data(c1_data[0][15:8])
    );
    
    pe u_pe_row0_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[2]),
        .in0_data(sys_arr_row0_data[23:16]),
        .in1_vld(sys_arr_col2_vld[0]),
        .in1_data(sys_arr_col2_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[2]),
        .out0_data(sys_arr_row1_data[23:16]),
        .out1_vld(sys_arr_col3_vld[0]),
        .out1_data(sys_arr_col3_data[7:0]),
        .pe_doing(pe_doing[0][2]),
        .c1_vld(c1_vld[0][2]),
        .c1_data(c1_data[0][23:16])
    );
    
    pe u_pe_row0_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[3]),
        .in0_data(sys_arr_row0_data[31:24]),
        .in1_vld(sys_arr_col3_vld[0]),
        .in1_data(sys_arr_col3_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[3]),
        .out0_data(sys_arr_row1_data[31:24]),
        .out1_vld(sys_arr_col4_vld[0]),
        .out1_data(sys_arr_col4_data[7:0]),
        .pe_doing(pe_doing[0][3]),
        .c1_vld(c1_vld[0][3]),
        .c1_data(c1_data[0][31:24])
    );
    
    pe u_pe_row0_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[4]),
        .in0_data(sys_arr_row0_data[39:32]),
        .in1_vld(sys_arr_col4_vld[0]),
        .in1_data(sys_arr_col4_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[4]),
        .out0_data(sys_arr_row1_data[39:32]),
        .out1_vld(sys_arr_col5_vld[0]),
        .out1_data(sys_arr_col5_data[7:0]),
        .pe_doing(pe_doing[0][4]),
        .c1_vld(c1_vld[0][4]),
        .c1_data(c1_data[0][39:32])
    );
    
    pe u_pe_row0_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[5]),
        .in0_data(sys_arr_row0_data[47:40]),
        .in1_vld(sys_arr_col5_vld[0]),
        .in1_data(sys_arr_col5_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[5]),
        .out0_data(sys_arr_row1_data[47:40]),
        .out1_vld(sys_arr_col6_vld[0]),
        .out1_data(sys_arr_col6_data[7:0]),
        .pe_doing(pe_doing[0][5]),
        .c1_vld(c1_vld[0][5]),
        .c1_data(c1_data[0][47:40])
    );
    
    pe u_pe_row0_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[6]),
        .in0_data(sys_arr_row0_data[55:48]),
        .in1_vld(sys_arr_col6_vld[0]),
        .in1_data(sys_arr_col6_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[6]),
        .out0_data(sys_arr_row1_data[55:48]),
        .out1_vld(sys_arr_col7_vld[0]),
        .out1_data(sys_arr_col7_data[7:0]),
        .pe_doing(pe_doing[0][6]),
        .c1_vld(c1_vld[0][6]),
        .c1_data(c1_data[0][55:48])
    );
    
    pe u_pe_row0_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[7]),
        .in0_data(sys_arr_row0_data[63:56]),
        .in1_vld(sys_arr_col7_vld[0]),
        .in1_data(sys_arr_col7_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[7]),
        .out0_data(sys_arr_row1_data[63:56]),
        .out1_vld(sys_arr_col8_vld[0]),
        .out1_data(sys_arr_col8_data[7:0]),
        .pe_doing(pe_doing[0][7]),
        .c1_vld(c1_vld[0][7]),
        .c1_data(c1_data[0][63:56])
    );
    
    pe u_pe_row0_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[8]),
        .in0_data(sys_arr_row0_data[71:64]),
        .in1_vld(sys_arr_col8_vld[0]),
        .in1_data(sys_arr_col8_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[8]),
        .out0_data(sys_arr_row1_data[71:64]),
        .out1_vld(sys_arr_col9_vld[0]),
        .out1_data(sys_arr_col9_data[7:0]),
        .pe_doing(pe_doing[0][8]),
        .c1_vld(c1_vld[0][8]),
        .c1_data(c1_data[0][71:64])
    );
    
    pe u_pe_row0_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[9]),
        .in0_data(sys_arr_row0_data[79:72]),
        .in1_vld(sys_arr_col9_vld[0]),
        .in1_data(sys_arr_col9_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[9]),
        .out0_data(sys_arr_row1_data[79:72]),
        .out1_vld(sys_arr_col10_vld[0]),
        .out1_data(sys_arr_col10_data[7:0]),
        .pe_doing(pe_doing[0][9]),
        .c1_vld(c1_vld[0][9]),
        .c1_data(c1_data[0][79:72])
    );
    
    pe u_pe_row0_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[10]),
        .in0_data(sys_arr_row0_data[87:80]),
        .in1_vld(sys_arr_col10_vld[0]),
        .in1_data(sys_arr_col10_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[10]),
        .out0_data(sys_arr_row1_data[87:80]),
        .out1_vld(sys_arr_col11_vld[0]),
        .out1_data(sys_arr_col11_data[7:0]),
        .pe_doing(pe_doing[0][10]),
        .c1_vld(c1_vld[0][10]),
        .c1_data(c1_data[0][87:80])
    );
    
    pe u_pe_row0_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[11]),
        .in0_data(sys_arr_row0_data[95:88]),
        .in1_vld(sys_arr_col11_vld[0]),
        .in1_data(sys_arr_col11_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[11]),
        .out0_data(sys_arr_row1_data[95:88]),
        .out1_vld(sys_arr_col12_vld[0]),
        .out1_data(sys_arr_col12_data[7:0]),
        .pe_doing(pe_doing[0][11]),
        .c1_vld(c1_vld[0][11]),
        .c1_data(c1_data[0][95:88])
    );
    
    pe u_pe_row0_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[12]),
        .in0_data(sys_arr_row0_data[103:96]),
        .in1_vld(sys_arr_col12_vld[0]),
        .in1_data(sys_arr_col12_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[12]),
        .out0_data(sys_arr_row1_data[103:96]),
        .out1_vld(sys_arr_col13_vld[0]),
        .out1_data(sys_arr_col13_data[7:0]),
        .pe_doing(pe_doing[0][12]),
        .c1_vld(c1_vld[0][12]),
        .c1_data(c1_data[0][103:96])
    );
    
    pe u_pe_row0_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[13]),
        .in0_data(sys_arr_row0_data[111:104]),
        .in1_vld(sys_arr_col13_vld[0]),
        .in1_data(sys_arr_col13_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[13]),
        .out0_data(sys_arr_row1_data[111:104]),
        .out1_vld(sys_arr_col14_vld[0]),
        .out1_data(sys_arr_col14_data[7:0]),
        .pe_doing(pe_doing[0][13]),
        .c1_vld(c1_vld[0][13]),
        .c1_data(c1_data[0][111:104])
    );
    
    pe u_pe_row0_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[14]),
        .in0_data(sys_arr_row0_data[119:112]),
        .in1_vld(sys_arr_col14_vld[0]),
        .in1_data(sys_arr_col14_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[14]),
        .out0_data(sys_arr_row1_data[119:112]),
        .out1_vld(sys_arr_col15_vld[0]),
        .out1_data(sys_arr_col15_data[7:0]),
        .pe_doing(pe_doing[0][14]),
        .c1_vld(c1_vld[0][14]),
        .c1_data(c1_data[0][119:112])
    );
    
    pe u_pe_row0_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row0_vld[15]),
        .in0_data(sys_arr_row0_data[127:120]),
        .in1_vld(sys_arr_col15_vld[0]),
        .in1_data(sys_arr_col15_data[7:0]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row1_vld[15]),
        .out0_data(sys_arr_row1_data[127:120]),
        .out1_vld(sys_arr_col16_vld[0]),
        .out1_data(sys_arr_col16_data[7:0]),
        .pe_doing(pe_doing[0][15]),
        .c1_vld(c1_vld[0][15]),
        .c1_data(c1_data[0][127:120])
    );
    
    pe u_pe_row1_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[0]),
        .in0_data(sys_arr_row1_data[7:0]),
        .in1_vld(sys_arr_col0_vld[1]),
        .in1_data(sys_arr_col0_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[0]),
        .out0_data(sys_arr_row2_data[7:0]),
        .out1_vld(sys_arr_col1_vld[1]),
        .out1_data(sys_arr_col1_data[15:8]),
        .pe_doing(pe_doing[1][0]),
        .c1_vld(c1_vld[1][0]),
        .c1_data(c1_data[1][7:0])
    );
    
    pe u_pe_row1_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[1]),
        .in0_data(sys_arr_row1_data[15:8]),
        .in1_vld(sys_arr_col1_vld[1]),
        .in1_data(sys_arr_col1_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[1]),
        .out0_data(sys_arr_row2_data[15:8]),
        .out1_vld(sys_arr_col2_vld[1]),
        .out1_data(sys_arr_col2_data[15:8]),
        .pe_doing(pe_doing[1][1]),
        .c1_vld(c1_vld[1][1]),
        .c1_data(c1_data[1][15:8])
    );
    
    pe u_pe_row1_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[2]),
        .in0_data(sys_arr_row1_data[23:16]),
        .in1_vld(sys_arr_col2_vld[1]),
        .in1_data(sys_arr_col2_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[2]),
        .out0_data(sys_arr_row2_data[23:16]),
        .out1_vld(sys_arr_col3_vld[1]),
        .out1_data(sys_arr_col3_data[15:8]),
        .pe_doing(pe_doing[1][2]),
        .c1_vld(c1_vld[1][2]),
        .c1_data(c1_data[1][23:16])
    );
    
    pe u_pe_row1_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[3]),
        .in0_data(sys_arr_row1_data[31:24]),
        .in1_vld(sys_arr_col3_vld[1]),
        .in1_data(sys_arr_col3_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[3]),
        .out0_data(sys_arr_row2_data[31:24]),
        .out1_vld(sys_arr_col4_vld[1]),
        .out1_data(sys_arr_col4_data[15:8]),
        .pe_doing(pe_doing[1][3]),
        .c1_vld(c1_vld[1][3]),
        .c1_data(c1_data[1][31:24])
    );
    
    pe u_pe_row1_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[4]),
        .in0_data(sys_arr_row1_data[39:32]),
        .in1_vld(sys_arr_col4_vld[1]),
        .in1_data(sys_arr_col4_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[4]),
        .out0_data(sys_arr_row2_data[39:32]),
        .out1_vld(sys_arr_col5_vld[1]),
        .out1_data(sys_arr_col5_data[15:8]),
        .pe_doing(pe_doing[1][4]),
        .c1_vld(c1_vld[1][4]),
        .c1_data(c1_data[1][39:32])
    );
    
    pe u_pe_row1_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[5]),
        .in0_data(sys_arr_row1_data[47:40]),
        .in1_vld(sys_arr_col5_vld[1]),
        .in1_data(sys_arr_col5_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[5]),
        .out0_data(sys_arr_row2_data[47:40]),
        .out1_vld(sys_arr_col6_vld[1]),
        .out1_data(sys_arr_col6_data[15:8]),
        .pe_doing(pe_doing[1][5]),
        .c1_vld(c1_vld[1][5]),
        .c1_data(c1_data[1][47:40])
    );
    
    pe u_pe_row1_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[6]),
        .in0_data(sys_arr_row1_data[55:48]),
        .in1_vld(sys_arr_col6_vld[1]),
        .in1_data(sys_arr_col6_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[6]),
        .out0_data(sys_arr_row2_data[55:48]),
        .out1_vld(sys_arr_col7_vld[1]),
        .out1_data(sys_arr_col7_data[15:8]),
        .pe_doing(pe_doing[1][6]),
        .c1_vld(c1_vld[1][6]),
        .c1_data(c1_data[1][55:48])
    );
    
    pe u_pe_row1_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[7]),
        .in0_data(sys_arr_row1_data[63:56]),
        .in1_vld(sys_arr_col7_vld[1]),
        .in1_data(sys_arr_col7_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[7]),
        .out0_data(sys_arr_row2_data[63:56]),
        .out1_vld(sys_arr_col8_vld[1]),
        .out1_data(sys_arr_col8_data[15:8]),
        .pe_doing(pe_doing[1][7]),
        .c1_vld(c1_vld[1][7]),
        .c1_data(c1_data[1][63:56])
    );
    
    pe u_pe_row1_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[8]),
        .in0_data(sys_arr_row1_data[71:64]),
        .in1_vld(sys_arr_col8_vld[1]),
        .in1_data(sys_arr_col8_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[8]),
        .out0_data(sys_arr_row2_data[71:64]),
        .out1_vld(sys_arr_col9_vld[1]),
        .out1_data(sys_arr_col9_data[15:8]),
        .pe_doing(pe_doing[1][8]),
        .c1_vld(c1_vld[1][8]),
        .c1_data(c1_data[1][71:64])
    );
    
    pe u_pe_row1_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[9]),
        .in0_data(sys_arr_row1_data[79:72]),
        .in1_vld(sys_arr_col9_vld[1]),
        .in1_data(sys_arr_col9_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[9]),
        .out0_data(sys_arr_row2_data[79:72]),
        .out1_vld(sys_arr_col10_vld[1]),
        .out1_data(sys_arr_col10_data[15:8]),
        .pe_doing(pe_doing[1][9]),
        .c1_vld(c1_vld[1][9]),
        .c1_data(c1_data[1][79:72])
    );
    
    pe u_pe_row1_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[10]),
        .in0_data(sys_arr_row1_data[87:80]),
        .in1_vld(sys_arr_col10_vld[1]),
        .in1_data(sys_arr_col10_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[10]),
        .out0_data(sys_arr_row2_data[87:80]),
        .out1_vld(sys_arr_col11_vld[1]),
        .out1_data(sys_arr_col11_data[15:8]),
        .pe_doing(pe_doing[1][10]),
        .c1_vld(c1_vld[1][10]),
        .c1_data(c1_data[1][87:80])
    );
    
    pe u_pe_row1_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[11]),
        .in0_data(sys_arr_row1_data[95:88]),
        .in1_vld(sys_arr_col11_vld[1]),
        .in1_data(sys_arr_col11_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[11]),
        .out0_data(sys_arr_row2_data[95:88]),
        .out1_vld(sys_arr_col12_vld[1]),
        .out1_data(sys_arr_col12_data[15:8]),
        .pe_doing(pe_doing[1][11]),
        .c1_vld(c1_vld[1][11]),
        .c1_data(c1_data[1][95:88])
    );
    
    pe u_pe_row1_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[12]),
        .in0_data(sys_arr_row1_data[103:96]),
        .in1_vld(sys_arr_col12_vld[1]),
        .in1_data(sys_arr_col12_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[12]),
        .out0_data(sys_arr_row2_data[103:96]),
        .out1_vld(sys_arr_col13_vld[1]),
        .out1_data(sys_arr_col13_data[15:8]),
        .pe_doing(pe_doing[1][12]),
        .c1_vld(c1_vld[1][12]),
        .c1_data(c1_data[1][103:96])
    );
    
    pe u_pe_row1_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[13]),
        .in0_data(sys_arr_row1_data[111:104]),
        .in1_vld(sys_arr_col13_vld[1]),
        .in1_data(sys_arr_col13_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[13]),
        .out0_data(sys_arr_row2_data[111:104]),
        .out1_vld(sys_arr_col14_vld[1]),
        .out1_data(sys_arr_col14_data[15:8]),
        .pe_doing(pe_doing[1][13]),
        .c1_vld(c1_vld[1][13]),
        .c1_data(c1_data[1][111:104])
    );
    
    pe u_pe_row1_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[14]),
        .in0_data(sys_arr_row1_data[119:112]),
        .in1_vld(sys_arr_col14_vld[1]),
        .in1_data(sys_arr_col14_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[14]),
        .out0_data(sys_arr_row2_data[119:112]),
        .out1_vld(sys_arr_col15_vld[1]),
        .out1_data(sys_arr_col15_data[15:8]),
        .pe_doing(pe_doing[1][14]),
        .c1_vld(c1_vld[1][14]),
        .c1_data(c1_data[1][119:112])
    );
    
    pe u_pe_row1_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row1_vld[15]),
        .in0_data(sys_arr_row1_data[127:120]),
        .in1_vld(sys_arr_col15_vld[1]),
        .in1_data(sys_arr_col15_data[15:8]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row2_vld[15]),
        .out0_data(sys_arr_row2_data[127:120]),
        .out1_vld(sys_arr_col16_vld[1]),
        .out1_data(sys_arr_col16_data[15:8]),
        .pe_doing(pe_doing[1][15]),
        .c1_vld(c1_vld[1][15]),
        .c1_data(c1_data[1][127:120])
    );
    
    pe u_pe_row2_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[0]),
        .in0_data(sys_arr_row2_data[7:0]),
        .in1_vld(sys_arr_col0_vld[2]),
        .in1_data(sys_arr_col0_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[0]),
        .out0_data(sys_arr_row3_data[7:0]),
        .out1_vld(sys_arr_col1_vld[2]),
        .out1_data(sys_arr_col1_data[23:16]),
        .pe_doing(pe_doing[2][0]),
        .c1_vld(c1_vld[2][0]),
        .c1_data(c1_data[2][7:0])
    );
    
    pe u_pe_row2_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[1]),
        .in0_data(sys_arr_row2_data[15:8]),
        .in1_vld(sys_arr_col1_vld[2]),
        .in1_data(sys_arr_col1_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[1]),
        .out0_data(sys_arr_row3_data[15:8]),
        .out1_vld(sys_arr_col2_vld[2]),
        .out1_data(sys_arr_col2_data[23:16]),
        .pe_doing(pe_doing[2][1]),
        .c1_vld(c1_vld[2][1]),
        .c1_data(c1_data[2][15:8])
    );
    
    pe u_pe_row2_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[2]),
        .in0_data(sys_arr_row2_data[23:16]),
        .in1_vld(sys_arr_col2_vld[2]),
        .in1_data(sys_arr_col2_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[2]),
        .out0_data(sys_arr_row3_data[23:16]),
        .out1_vld(sys_arr_col3_vld[2]),
        .out1_data(sys_arr_col3_data[23:16]),
        .pe_doing(pe_doing[2][2]),
        .c1_vld(c1_vld[2][2]),
        .c1_data(c1_data[2][23:16])
    );
    
    pe u_pe_row2_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[3]),
        .in0_data(sys_arr_row2_data[31:24]),
        .in1_vld(sys_arr_col3_vld[2]),
        .in1_data(sys_arr_col3_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[3]),
        .out0_data(sys_arr_row3_data[31:24]),
        .out1_vld(sys_arr_col4_vld[2]),
        .out1_data(sys_arr_col4_data[23:16]),
        .pe_doing(pe_doing[2][3]),
        .c1_vld(c1_vld[2][3]),
        .c1_data(c1_data[2][31:24])
    );
    
    pe u_pe_row2_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[4]),
        .in0_data(sys_arr_row2_data[39:32]),
        .in1_vld(sys_arr_col4_vld[2]),
        .in1_data(sys_arr_col4_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[4]),
        .out0_data(sys_arr_row3_data[39:32]),
        .out1_vld(sys_arr_col5_vld[2]),
        .out1_data(sys_arr_col5_data[23:16]),
        .pe_doing(pe_doing[2][4]),
        .c1_vld(c1_vld[2][4]),
        .c1_data(c1_data[2][39:32])
    );
    
    pe u_pe_row2_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[5]),
        .in0_data(sys_arr_row2_data[47:40]),
        .in1_vld(sys_arr_col5_vld[2]),
        .in1_data(sys_arr_col5_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[5]),
        .out0_data(sys_arr_row3_data[47:40]),
        .out1_vld(sys_arr_col6_vld[2]),
        .out1_data(sys_arr_col6_data[23:16]),
        .pe_doing(pe_doing[2][5]),
        .c1_vld(c1_vld[2][5]),
        .c1_data(c1_data[2][47:40])
    );
    
    pe u_pe_row2_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[6]),
        .in0_data(sys_arr_row2_data[55:48]),
        .in1_vld(sys_arr_col6_vld[2]),
        .in1_data(sys_arr_col6_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[6]),
        .out0_data(sys_arr_row3_data[55:48]),
        .out1_vld(sys_arr_col7_vld[2]),
        .out1_data(sys_arr_col7_data[23:16]),
        .pe_doing(pe_doing[2][6]),
        .c1_vld(c1_vld[2][6]),
        .c1_data(c1_data[2][55:48])
    );
    
    pe u_pe_row2_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[7]),
        .in0_data(sys_arr_row2_data[63:56]),
        .in1_vld(sys_arr_col7_vld[2]),
        .in1_data(sys_arr_col7_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[7]),
        .out0_data(sys_arr_row3_data[63:56]),
        .out1_vld(sys_arr_col8_vld[2]),
        .out1_data(sys_arr_col8_data[23:16]),
        .pe_doing(pe_doing[2][7]),
        .c1_vld(c1_vld[2][7]),
        .c1_data(c1_data[2][63:56])
    );
    
    pe u_pe_row2_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[8]),
        .in0_data(sys_arr_row2_data[71:64]),
        .in1_vld(sys_arr_col8_vld[2]),
        .in1_data(sys_arr_col8_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[8]),
        .out0_data(sys_arr_row3_data[71:64]),
        .out1_vld(sys_arr_col9_vld[2]),
        .out1_data(sys_arr_col9_data[23:16]),
        .pe_doing(pe_doing[2][8]),
        .c1_vld(c1_vld[2][8]),
        .c1_data(c1_data[2][71:64])
    );
    
    pe u_pe_row2_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[9]),
        .in0_data(sys_arr_row2_data[79:72]),
        .in1_vld(sys_arr_col9_vld[2]),
        .in1_data(sys_arr_col9_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[9]),
        .out0_data(sys_arr_row3_data[79:72]),
        .out1_vld(sys_arr_col10_vld[2]),
        .out1_data(sys_arr_col10_data[23:16]),
        .pe_doing(pe_doing[2][9]),
        .c1_vld(c1_vld[2][9]),
        .c1_data(c1_data[2][79:72])
    );
    
    pe u_pe_row2_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[10]),
        .in0_data(sys_arr_row2_data[87:80]),
        .in1_vld(sys_arr_col10_vld[2]),
        .in1_data(sys_arr_col10_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[10]),
        .out0_data(sys_arr_row3_data[87:80]),
        .out1_vld(sys_arr_col11_vld[2]),
        .out1_data(sys_arr_col11_data[23:16]),
        .pe_doing(pe_doing[2][10]),
        .c1_vld(c1_vld[2][10]),
        .c1_data(c1_data[2][87:80])
    );
    
    pe u_pe_row2_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[11]),
        .in0_data(sys_arr_row2_data[95:88]),
        .in1_vld(sys_arr_col11_vld[2]),
        .in1_data(sys_arr_col11_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[11]),
        .out0_data(sys_arr_row3_data[95:88]),
        .out1_vld(sys_arr_col12_vld[2]),
        .out1_data(sys_arr_col12_data[23:16]),
        .pe_doing(pe_doing[2][11]),
        .c1_vld(c1_vld[2][11]),
        .c1_data(c1_data[2][95:88])
    );
    
    pe u_pe_row2_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[12]),
        .in0_data(sys_arr_row2_data[103:96]),
        .in1_vld(sys_arr_col12_vld[2]),
        .in1_data(sys_arr_col12_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[12]),
        .out0_data(sys_arr_row3_data[103:96]),
        .out1_vld(sys_arr_col13_vld[2]),
        .out1_data(sys_arr_col13_data[23:16]),
        .pe_doing(pe_doing[2][12]),
        .c1_vld(c1_vld[2][12]),
        .c1_data(c1_data[2][103:96])
    );
    
    pe u_pe_row2_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[13]),
        .in0_data(sys_arr_row2_data[111:104]),
        .in1_vld(sys_arr_col13_vld[2]),
        .in1_data(sys_arr_col13_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[13]),
        .out0_data(sys_arr_row3_data[111:104]),
        .out1_vld(sys_arr_col14_vld[2]),
        .out1_data(sys_arr_col14_data[23:16]),
        .pe_doing(pe_doing[2][13]),
        .c1_vld(c1_vld[2][13]),
        .c1_data(c1_data[2][111:104])
    );
    
    pe u_pe_row2_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[14]),
        .in0_data(sys_arr_row2_data[119:112]),
        .in1_vld(sys_arr_col14_vld[2]),
        .in1_data(sys_arr_col14_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[14]),
        .out0_data(sys_arr_row3_data[119:112]),
        .out1_vld(sys_arr_col15_vld[2]),
        .out1_data(sys_arr_col15_data[23:16]),
        .pe_doing(pe_doing[2][14]),
        .c1_vld(c1_vld[2][14]),
        .c1_data(c1_data[2][119:112])
    );
    
    pe u_pe_row2_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row2_vld[15]),
        .in0_data(sys_arr_row2_data[127:120]),
        .in1_vld(sys_arr_col15_vld[2]),
        .in1_data(sys_arr_col15_data[23:16]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row3_vld[15]),
        .out0_data(sys_arr_row3_data[127:120]),
        .out1_vld(sys_arr_col16_vld[2]),
        .out1_data(sys_arr_col16_data[23:16]),
        .pe_doing(pe_doing[2][15]),
        .c1_vld(c1_vld[2][15]),
        .c1_data(c1_data[2][127:120])
    );
    
    pe u_pe_row3_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[0]),
        .in0_data(sys_arr_row3_data[7:0]),
        .in1_vld(sys_arr_col0_vld[3]),
        .in1_data(sys_arr_col0_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[0]),
        .out0_data(sys_arr_row4_data[7:0]),
        .out1_vld(sys_arr_col1_vld[3]),
        .out1_data(sys_arr_col1_data[31:24]),
        .pe_doing(pe_doing[3][0]),
        .c1_vld(c1_vld[3][0]),
        .c1_data(c1_data[3][7:0])
    );
    
    pe u_pe_row3_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[1]),
        .in0_data(sys_arr_row3_data[15:8]),
        .in1_vld(sys_arr_col1_vld[3]),
        .in1_data(sys_arr_col1_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[1]),
        .out0_data(sys_arr_row4_data[15:8]),
        .out1_vld(sys_arr_col2_vld[3]),
        .out1_data(sys_arr_col2_data[31:24]),
        .pe_doing(pe_doing[3][1]),
        .c1_vld(c1_vld[3][1]),
        .c1_data(c1_data[3][15:8])
    );
    
    pe u_pe_row3_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[2]),
        .in0_data(sys_arr_row3_data[23:16]),
        .in1_vld(sys_arr_col2_vld[3]),
        .in1_data(sys_arr_col2_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[2]),
        .out0_data(sys_arr_row4_data[23:16]),
        .out1_vld(sys_arr_col3_vld[3]),
        .out1_data(sys_arr_col3_data[31:24]),
        .pe_doing(pe_doing[3][2]),
        .c1_vld(c1_vld[3][2]),
        .c1_data(c1_data[3][23:16])
    );
    
    pe u_pe_row3_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[3]),
        .in0_data(sys_arr_row3_data[31:24]),
        .in1_vld(sys_arr_col3_vld[3]),
        .in1_data(sys_arr_col3_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[3]),
        .out0_data(sys_arr_row4_data[31:24]),
        .out1_vld(sys_arr_col4_vld[3]),
        .out1_data(sys_arr_col4_data[31:24]),
        .pe_doing(pe_doing[3][3]),
        .c1_vld(c1_vld[3][3]),
        .c1_data(c1_data[3][31:24])
    );
    
    pe u_pe_row3_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[4]),
        .in0_data(sys_arr_row3_data[39:32]),
        .in1_vld(sys_arr_col4_vld[3]),
        .in1_data(sys_arr_col4_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[4]),
        .out0_data(sys_arr_row4_data[39:32]),
        .out1_vld(sys_arr_col5_vld[3]),
        .out1_data(sys_arr_col5_data[31:24]),
        .pe_doing(pe_doing[3][4]),
        .c1_vld(c1_vld[3][4]),
        .c1_data(c1_data[3][39:32])
    );
    
    pe u_pe_row3_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[5]),
        .in0_data(sys_arr_row3_data[47:40]),
        .in1_vld(sys_arr_col5_vld[3]),
        .in1_data(sys_arr_col5_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[5]),
        .out0_data(sys_arr_row4_data[47:40]),
        .out1_vld(sys_arr_col6_vld[3]),
        .out1_data(sys_arr_col6_data[31:24]),
        .pe_doing(pe_doing[3][5]),
        .c1_vld(c1_vld[3][5]),
        .c1_data(c1_data[3][47:40])
    );
    
    pe u_pe_row3_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[6]),
        .in0_data(sys_arr_row3_data[55:48]),
        .in1_vld(sys_arr_col6_vld[3]),
        .in1_data(sys_arr_col6_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[6]),
        .out0_data(sys_arr_row4_data[55:48]),
        .out1_vld(sys_arr_col7_vld[3]),
        .out1_data(sys_arr_col7_data[31:24]),
        .pe_doing(pe_doing[3][6]),
        .c1_vld(c1_vld[3][6]),
        .c1_data(c1_data[3][55:48])
    );
    
    pe u_pe_row3_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[7]),
        .in0_data(sys_arr_row3_data[63:56]),
        .in1_vld(sys_arr_col7_vld[3]),
        .in1_data(sys_arr_col7_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[7]),
        .out0_data(sys_arr_row4_data[63:56]),
        .out1_vld(sys_arr_col8_vld[3]),
        .out1_data(sys_arr_col8_data[31:24]),
        .pe_doing(pe_doing[3][7]),
        .c1_vld(c1_vld[3][7]),
        .c1_data(c1_data[3][63:56])
    );
    
    pe u_pe_row3_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[8]),
        .in0_data(sys_arr_row3_data[71:64]),
        .in1_vld(sys_arr_col8_vld[3]),
        .in1_data(sys_arr_col8_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[8]),
        .out0_data(sys_arr_row4_data[71:64]),
        .out1_vld(sys_arr_col9_vld[3]),
        .out1_data(sys_arr_col9_data[31:24]),
        .pe_doing(pe_doing[3][8]),
        .c1_vld(c1_vld[3][8]),
        .c1_data(c1_data[3][71:64])
    );
    
    pe u_pe_row3_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[9]),
        .in0_data(sys_arr_row3_data[79:72]),
        .in1_vld(sys_arr_col9_vld[3]),
        .in1_data(sys_arr_col9_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[9]),
        .out0_data(sys_arr_row4_data[79:72]),
        .out1_vld(sys_arr_col10_vld[3]),
        .out1_data(sys_arr_col10_data[31:24]),
        .pe_doing(pe_doing[3][9]),
        .c1_vld(c1_vld[3][9]),
        .c1_data(c1_data[3][79:72])
    );
    
    pe u_pe_row3_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[10]),
        .in0_data(sys_arr_row3_data[87:80]),
        .in1_vld(sys_arr_col10_vld[3]),
        .in1_data(sys_arr_col10_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[10]),
        .out0_data(sys_arr_row4_data[87:80]),
        .out1_vld(sys_arr_col11_vld[3]),
        .out1_data(sys_arr_col11_data[31:24]),
        .pe_doing(pe_doing[3][10]),
        .c1_vld(c1_vld[3][10]),
        .c1_data(c1_data[3][87:80])
    );
    
    pe u_pe_row3_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[11]),
        .in0_data(sys_arr_row3_data[95:88]),
        .in1_vld(sys_arr_col11_vld[3]),
        .in1_data(sys_arr_col11_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[11]),
        .out0_data(sys_arr_row4_data[95:88]),
        .out1_vld(sys_arr_col12_vld[3]),
        .out1_data(sys_arr_col12_data[31:24]),
        .pe_doing(pe_doing[3][11]),
        .c1_vld(c1_vld[3][11]),
        .c1_data(c1_data[3][95:88])
    );
    
    pe u_pe_row3_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[12]),
        .in0_data(sys_arr_row3_data[103:96]),
        .in1_vld(sys_arr_col12_vld[3]),
        .in1_data(sys_arr_col12_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[12]),
        .out0_data(sys_arr_row4_data[103:96]),
        .out1_vld(sys_arr_col13_vld[3]),
        .out1_data(sys_arr_col13_data[31:24]),
        .pe_doing(pe_doing[3][12]),
        .c1_vld(c1_vld[3][12]),
        .c1_data(c1_data[3][103:96])
    );
    
    pe u_pe_row3_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[13]),
        .in0_data(sys_arr_row3_data[111:104]),
        .in1_vld(sys_arr_col13_vld[3]),
        .in1_data(sys_arr_col13_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[13]),
        .out0_data(sys_arr_row4_data[111:104]),
        .out1_vld(sys_arr_col14_vld[3]),
        .out1_data(sys_arr_col14_data[31:24]),
        .pe_doing(pe_doing[3][13]),
        .c1_vld(c1_vld[3][13]),
        .c1_data(c1_data[3][111:104])
    );
    
    pe u_pe_row3_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[14]),
        .in0_data(sys_arr_row3_data[119:112]),
        .in1_vld(sys_arr_col14_vld[3]),
        .in1_data(sys_arr_col14_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[14]),
        .out0_data(sys_arr_row4_data[119:112]),
        .out1_vld(sys_arr_col15_vld[3]),
        .out1_data(sys_arr_col15_data[31:24]),
        .pe_doing(pe_doing[3][14]),
        .c1_vld(c1_vld[3][14]),
        .c1_data(c1_data[3][119:112])
    );
    
    pe u_pe_row3_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row3_vld[15]),
        .in0_data(sys_arr_row3_data[127:120]),
        .in1_vld(sys_arr_col15_vld[3]),
        .in1_data(sys_arr_col15_data[31:24]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row4_vld[15]),
        .out0_data(sys_arr_row4_data[127:120]),
        .out1_vld(sys_arr_col16_vld[3]),
        .out1_data(sys_arr_col16_data[31:24]),
        .pe_doing(pe_doing[3][15]),
        .c1_vld(c1_vld[3][15]),
        .c1_data(c1_data[3][127:120])
    );
    
    pe u_pe_row4_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[0]),
        .in0_data(sys_arr_row4_data[7:0]),
        .in1_vld(sys_arr_col0_vld[4]),
        .in1_data(sys_arr_col0_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[0]),
        .out0_data(sys_arr_row5_data[7:0]),
        .out1_vld(sys_arr_col1_vld[4]),
        .out1_data(sys_arr_col1_data[39:32]),
        .pe_doing(pe_doing[4][0]),
        .c1_vld(c1_vld[4][0]),
        .c1_data(c1_data[4][7:0])
    );
    
    pe u_pe_row4_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[1]),
        .in0_data(sys_arr_row4_data[15:8]),
        .in1_vld(sys_arr_col1_vld[4]),
        .in1_data(sys_arr_col1_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[1]),
        .out0_data(sys_arr_row5_data[15:8]),
        .out1_vld(sys_arr_col2_vld[4]),
        .out1_data(sys_arr_col2_data[39:32]),
        .pe_doing(pe_doing[4][1]),
        .c1_vld(c1_vld[4][1]),
        .c1_data(c1_data[4][15:8])
    );
    
    pe u_pe_row4_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[2]),
        .in0_data(sys_arr_row4_data[23:16]),
        .in1_vld(sys_arr_col2_vld[4]),
        .in1_data(sys_arr_col2_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[2]),
        .out0_data(sys_arr_row5_data[23:16]),
        .out1_vld(sys_arr_col3_vld[4]),
        .out1_data(sys_arr_col3_data[39:32]),
        .pe_doing(pe_doing[4][2]),
        .c1_vld(c1_vld[4][2]),
        .c1_data(c1_data[4][23:16])
    );
    
    pe u_pe_row4_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[3]),
        .in0_data(sys_arr_row4_data[31:24]),
        .in1_vld(sys_arr_col3_vld[4]),
        .in1_data(sys_arr_col3_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[3]),
        .out0_data(sys_arr_row5_data[31:24]),
        .out1_vld(sys_arr_col4_vld[4]),
        .out1_data(sys_arr_col4_data[39:32]),
        .pe_doing(pe_doing[4][3]),
        .c1_vld(c1_vld[4][3]),
        .c1_data(c1_data[4][31:24])
    );
    
    pe u_pe_row4_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[4]),
        .in0_data(sys_arr_row4_data[39:32]),
        .in1_vld(sys_arr_col4_vld[4]),
        .in1_data(sys_arr_col4_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[4]),
        .out0_data(sys_arr_row5_data[39:32]),
        .out1_vld(sys_arr_col5_vld[4]),
        .out1_data(sys_arr_col5_data[39:32]),
        .pe_doing(pe_doing[4][4]),
        .c1_vld(c1_vld[4][4]),
        .c1_data(c1_data[4][39:32])
    );
    
    pe u_pe_row4_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[5]),
        .in0_data(sys_arr_row4_data[47:40]),
        .in1_vld(sys_arr_col5_vld[4]),
        .in1_data(sys_arr_col5_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[5]),
        .out0_data(sys_arr_row5_data[47:40]),
        .out1_vld(sys_arr_col6_vld[4]),
        .out1_data(sys_arr_col6_data[39:32]),
        .pe_doing(pe_doing[4][5]),
        .c1_vld(c1_vld[4][5]),
        .c1_data(c1_data[4][47:40])
    );
    
    pe u_pe_row4_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[6]),
        .in0_data(sys_arr_row4_data[55:48]),
        .in1_vld(sys_arr_col6_vld[4]),
        .in1_data(sys_arr_col6_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[6]),
        .out0_data(sys_arr_row5_data[55:48]),
        .out1_vld(sys_arr_col7_vld[4]),
        .out1_data(sys_arr_col7_data[39:32]),
        .pe_doing(pe_doing[4][6]),
        .c1_vld(c1_vld[4][6]),
        .c1_data(c1_data[4][55:48])
    );
    
    pe u_pe_row4_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[7]),
        .in0_data(sys_arr_row4_data[63:56]),
        .in1_vld(sys_arr_col7_vld[4]),
        .in1_data(sys_arr_col7_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[7]),
        .out0_data(sys_arr_row5_data[63:56]),
        .out1_vld(sys_arr_col8_vld[4]),
        .out1_data(sys_arr_col8_data[39:32]),
        .pe_doing(pe_doing[4][7]),
        .c1_vld(c1_vld[4][7]),
        .c1_data(c1_data[4][63:56])
    );
    
    pe u_pe_row4_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[8]),
        .in0_data(sys_arr_row4_data[71:64]),
        .in1_vld(sys_arr_col8_vld[4]),
        .in1_data(sys_arr_col8_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[8]),
        .out0_data(sys_arr_row5_data[71:64]),
        .out1_vld(sys_arr_col9_vld[4]),
        .out1_data(sys_arr_col9_data[39:32]),
        .pe_doing(pe_doing[4][8]),
        .c1_vld(c1_vld[4][8]),
        .c1_data(c1_data[4][71:64])
    );
    
    pe u_pe_row4_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[9]),
        .in0_data(sys_arr_row4_data[79:72]),
        .in1_vld(sys_arr_col9_vld[4]),
        .in1_data(sys_arr_col9_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[9]),
        .out0_data(sys_arr_row5_data[79:72]),
        .out1_vld(sys_arr_col10_vld[4]),
        .out1_data(sys_arr_col10_data[39:32]),
        .pe_doing(pe_doing[4][9]),
        .c1_vld(c1_vld[4][9]),
        .c1_data(c1_data[4][79:72])
    );
    
    pe u_pe_row4_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[10]),
        .in0_data(sys_arr_row4_data[87:80]),
        .in1_vld(sys_arr_col10_vld[4]),
        .in1_data(sys_arr_col10_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[10]),
        .out0_data(sys_arr_row5_data[87:80]),
        .out1_vld(sys_arr_col11_vld[4]),
        .out1_data(sys_arr_col11_data[39:32]),
        .pe_doing(pe_doing[4][10]),
        .c1_vld(c1_vld[4][10]),
        .c1_data(c1_data[4][87:80])
    );
    
    pe u_pe_row4_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[11]),
        .in0_data(sys_arr_row4_data[95:88]),
        .in1_vld(sys_arr_col11_vld[4]),
        .in1_data(sys_arr_col11_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[11]),
        .out0_data(sys_arr_row5_data[95:88]),
        .out1_vld(sys_arr_col12_vld[4]),
        .out1_data(sys_arr_col12_data[39:32]),
        .pe_doing(pe_doing[4][11]),
        .c1_vld(c1_vld[4][11]),
        .c1_data(c1_data[4][95:88])
    );
    
    pe u_pe_row4_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[12]),
        .in0_data(sys_arr_row4_data[103:96]),
        .in1_vld(sys_arr_col12_vld[4]),
        .in1_data(sys_arr_col12_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[12]),
        .out0_data(sys_arr_row5_data[103:96]),
        .out1_vld(sys_arr_col13_vld[4]),
        .out1_data(sys_arr_col13_data[39:32]),
        .pe_doing(pe_doing[4][12]),
        .c1_vld(c1_vld[4][12]),
        .c1_data(c1_data[4][103:96])
    );
    
    pe u_pe_row4_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[13]),
        .in0_data(sys_arr_row4_data[111:104]),
        .in1_vld(sys_arr_col13_vld[4]),
        .in1_data(sys_arr_col13_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[13]),
        .out0_data(sys_arr_row5_data[111:104]),
        .out1_vld(sys_arr_col14_vld[4]),
        .out1_data(sys_arr_col14_data[39:32]),
        .pe_doing(pe_doing[4][13]),
        .c1_vld(c1_vld[4][13]),
        .c1_data(c1_data[4][111:104])
    );
    
    pe u_pe_row4_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[14]),
        .in0_data(sys_arr_row4_data[119:112]),
        .in1_vld(sys_arr_col14_vld[4]),
        .in1_data(sys_arr_col14_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[14]),
        .out0_data(sys_arr_row5_data[119:112]),
        .out1_vld(sys_arr_col15_vld[4]),
        .out1_data(sys_arr_col15_data[39:32]),
        .pe_doing(pe_doing[4][14]),
        .c1_vld(c1_vld[4][14]),
        .c1_data(c1_data[4][119:112])
    );
    
    pe u_pe_row4_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row4_vld[15]),
        .in0_data(sys_arr_row4_data[127:120]),
        .in1_vld(sys_arr_col15_vld[4]),
        .in1_data(sys_arr_col15_data[39:32]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row5_vld[15]),
        .out0_data(sys_arr_row5_data[127:120]),
        .out1_vld(sys_arr_col16_vld[4]),
        .out1_data(sys_arr_col16_data[39:32]),
        .pe_doing(pe_doing[4][15]),
        .c1_vld(c1_vld[4][15]),
        .c1_data(c1_data[4][127:120])
    );
    
    pe u_pe_row5_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[0]),
        .in0_data(sys_arr_row5_data[7:0]),
        .in1_vld(sys_arr_col0_vld[5]),
        .in1_data(sys_arr_col0_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[0]),
        .out0_data(sys_arr_row6_data[7:0]),
        .out1_vld(sys_arr_col1_vld[5]),
        .out1_data(sys_arr_col1_data[47:40]),
        .pe_doing(pe_doing[5][0]),
        .c1_vld(c1_vld[5][0]),
        .c1_data(c1_data[5][7:0])
    );
    
    pe u_pe_row5_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[1]),
        .in0_data(sys_arr_row5_data[15:8]),
        .in1_vld(sys_arr_col1_vld[5]),
        .in1_data(sys_arr_col1_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[1]),
        .out0_data(sys_arr_row6_data[15:8]),
        .out1_vld(sys_arr_col2_vld[5]),
        .out1_data(sys_arr_col2_data[47:40]),
        .pe_doing(pe_doing[5][1]),
        .c1_vld(c1_vld[5][1]),
        .c1_data(c1_data[5][15:8])
    );
    
    pe u_pe_row5_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[2]),
        .in0_data(sys_arr_row5_data[23:16]),
        .in1_vld(sys_arr_col2_vld[5]),
        .in1_data(sys_arr_col2_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[2]),
        .out0_data(sys_arr_row6_data[23:16]),
        .out1_vld(sys_arr_col3_vld[5]),
        .out1_data(sys_arr_col3_data[47:40]),
        .pe_doing(pe_doing[5][2]),
        .c1_vld(c1_vld[5][2]),
        .c1_data(c1_data[5][23:16])
    );
    
    pe u_pe_row5_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[3]),
        .in0_data(sys_arr_row5_data[31:24]),
        .in1_vld(sys_arr_col3_vld[5]),
        .in1_data(sys_arr_col3_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[3]),
        .out0_data(sys_arr_row6_data[31:24]),
        .out1_vld(sys_arr_col4_vld[5]),
        .out1_data(sys_arr_col4_data[47:40]),
        .pe_doing(pe_doing[5][3]),
        .c1_vld(c1_vld[5][3]),
        .c1_data(c1_data[5][31:24])
    );
    
    pe u_pe_row5_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[4]),
        .in0_data(sys_arr_row5_data[39:32]),
        .in1_vld(sys_arr_col4_vld[5]),
        .in1_data(sys_arr_col4_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[4]),
        .out0_data(sys_arr_row6_data[39:32]),
        .out1_vld(sys_arr_col5_vld[5]),
        .out1_data(sys_arr_col5_data[47:40]),
        .pe_doing(pe_doing[5][4]),
        .c1_vld(c1_vld[5][4]),
        .c1_data(c1_data[5][39:32])
    );
    
    pe u_pe_row5_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[5]),
        .in0_data(sys_arr_row5_data[47:40]),
        .in1_vld(sys_arr_col5_vld[5]),
        .in1_data(sys_arr_col5_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[5]),
        .out0_data(sys_arr_row6_data[47:40]),
        .out1_vld(sys_arr_col6_vld[5]),
        .out1_data(sys_arr_col6_data[47:40]),
        .pe_doing(pe_doing[5][5]),
        .c1_vld(c1_vld[5][5]),
        .c1_data(c1_data[5][47:40])
    );
    
    pe u_pe_row5_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[6]),
        .in0_data(sys_arr_row5_data[55:48]),
        .in1_vld(sys_arr_col6_vld[5]),
        .in1_data(sys_arr_col6_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[6]),
        .out0_data(sys_arr_row6_data[55:48]),
        .out1_vld(sys_arr_col7_vld[5]),
        .out1_data(sys_arr_col7_data[47:40]),
        .pe_doing(pe_doing[5][6]),
        .c1_vld(c1_vld[5][6]),
        .c1_data(c1_data[5][55:48])
    );
    
    pe u_pe_row5_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[7]),
        .in0_data(sys_arr_row5_data[63:56]),
        .in1_vld(sys_arr_col7_vld[5]),
        .in1_data(sys_arr_col7_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[7]),
        .out0_data(sys_arr_row6_data[63:56]),
        .out1_vld(sys_arr_col8_vld[5]),
        .out1_data(sys_arr_col8_data[47:40]),
        .pe_doing(pe_doing[5][7]),
        .c1_vld(c1_vld[5][7]),
        .c1_data(c1_data[5][63:56])
    );
    
    pe u_pe_row5_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[8]),
        .in0_data(sys_arr_row5_data[71:64]),
        .in1_vld(sys_arr_col8_vld[5]),
        .in1_data(sys_arr_col8_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[8]),
        .out0_data(sys_arr_row6_data[71:64]),
        .out1_vld(sys_arr_col9_vld[5]),
        .out1_data(sys_arr_col9_data[47:40]),
        .pe_doing(pe_doing[5][8]),
        .c1_vld(c1_vld[5][8]),
        .c1_data(c1_data[5][71:64])
    );
    
    pe u_pe_row5_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[9]),
        .in0_data(sys_arr_row5_data[79:72]),
        .in1_vld(sys_arr_col9_vld[5]),
        .in1_data(sys_arr_col9_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[9]),
        .out0_data(sys_arr_row6_data[79:72]),
        .out1_vld(sys_arr_col10_vld[5]),
        .out1_data(sys_arr_col10_data[47:40]),
        .pe_doing(pe_doing[5][9]),
        .c1_vld(c1_vld[5][9]),
        .c1_data(c1_data[5][79:72])
    );
    
    pe u_pe_row5_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[10]),
        .in0_data(sys_arr_row5_data[87:80]),
        .in1_vld(sys_arr_col10_vld[5]),
        .in1_data(sys_arr_col10_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[10]),
        .out0_data(sys_arr_row6_data[87:80]),
        .out1_vld(sys_arr_col11_vld[5]),
        .out1_data(sys_arr_col11_data[47:40]),
        .pe_doing(pe_doing[5][10]),
        .c1_vld(c1_vld[5][10]),
        .c1_data(c1_data[5][87:80])
    );
    
    pe u_pe_row5_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[11]),
        .in0_data(sys_arr_row5_data[95:88]),
        .in1_vld(sys_arr_col11_vld[5]),
        .in1_data(sys_arr_col11_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[11]),
        .out0_data(sys_arr_row6_data[95:88]),
        .out1_vld(sys_arr_col12_vld[5]),
        .out1_data(sys_arr_col12_data[47:40]),
        .pe_doing(pe_doing[5][11]),
        .c1_vld(c1_vld[5][11]),
        .c1_data(c1_data[5][95:88])
    );
    
    pe u_pe_row5_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[12]),
        .in0_data(sys_arr_row5_data[103:96]),
        .in1_vld(sys_arr_col12_vld[5]),
        .in1_data(sys_arr_col12_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[12]),
        .out0_data(sys_arr_row6_data[103:96]),
        .out1_vld(sys_arr_col13_vld[5]),
        .out1_data(sys_arr_col13_data[47:40]),
        .pe_doing(pe_doing[5][12]),
        .c1_vld(c1_vld[5][12]),
        .c1_data(c1_data[5][103:96])
    );
    
    pe u_pe_row5_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[13]),
        .in0_data(sys_arr_row5_data[111:104]),
        .in1_vld(sys_arr_col13_vld[5]),
        .in1_data(sys_arr_col13_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[13]),
        .out0_data(sys_arr_row6_data[111:104]),
        .out1_vld(sys_arr_col14_vld[5]),
        .out1_data(sys_arr_col14_data[47:40]),
        .pe_doing(pe_doing[5][13]),
        .c1_vld(c1_vld[5][13]),
        .c1_data(c1_data[5][111:104])
    );
    
    pe u_pe_row5_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[14]),
        .in0_data(sys_arr_row5_data[119:112]),
        .in1_vld(sys_arr_col14_vld[5]),
        .in1_data(sys_arr_col14_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[14]),
        .out0_data(sys_arr_row6_data[119:112]),
        .out1_vld(sys_arr_col15_vld[5]),
        .out1_data(sys_arr_col15_data[47:40]),
        .pe_doing(pe_doing[5][14]),
        .c1_vld(c1_vld[5][14]),
        .c1_data(c1_data[5][119:112])
    );
    
    pe u_pe_row5_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row5_vld[15]),
        .in0_data(sys_arr_row5_data[127:120]),
        .in1_vld(sys_arr_col15_vld[5]),
        .in1_data(sys_arr_col15_data[47:40]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row6_vld[15]),
        .out0_data(sys_arr_row6_data[127:120]),
        .out1_vld(sys_arr_col16_vld[5]),
        .out1_data(sys_arr_col16_data[47:40]),
        .pe_doing(pe_doing[5][15]),
        .c1_vld(c1_vld[5][15]),
        .c1_data(c1_data[5][127:120])
    );
    
    pe u_pe_row6_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[0]),
        .in0_data(sys_arr_row6_data[7:0]),
        .in1_vld(sys_arr_col0_vld[6]),
        .in1_data(sys_arr_col0_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[0]),
        .out0_data(sys_arr_row7_data[7:0]),
        .out1_vld(sys_arr_col1_vld[6]),
        .out1_data(sys_arr_col1_data[55:48]),
        .pe_doing(pe_doing[6][0]),
        .c1_vld(c1_vld[6][0]),
        .c1_data(c1_data[6][7:0])
    );
    
    pe u_pe_row6_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[1]),
        .in0_data(sys_arr_row6_data[15:8]),
        .in1_vld(sys_arr_col1_vld[6]),
        .in1_data(sys_arr_col1_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[1]),
        .out0_data(sys_arr_row7_data[15:8]),
        .out1_vld(sys_arr_col2_vld[6]),
        .out1_data(sys_arr_col2_data[55:48]),
        .pe_doing(pe_doing[6][1]),
        .c1_vld(c1_vld[6][1]),
        .c1_data(c1_data[6][15:8])
    );
    
    pe u_pe_row6_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[2]),
        .in0_data(sys_arr_row6_data[23:16]),
        .in1_vld(sys_arr_col2_vld[6]),
        .in1_data(sys_arr_col2_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[2]),
        .out0_data(sys_arr_row7_data[23:16]),
        .out1_vld(sys_arr_col3_vld[6]),
        .out1_data(sys_arr_col3_data[55:48]),
        .pe_doing(pe_doing[6][2]),
        .c1_vld(c1_vld[6][2]),
        .c1_data(c1_data[6][23:16])
    );
    
    pe u_pe_row6_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[3]),
        .in0_data(sys_arr_row6_data[31:24]),
        .in1_vld(sys_arr_col3_vld[6]),
        .in1_data(sys_arr_col3_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[3]),
        .out0_data(sys_arr_row7_data[31:24]),
        .out1_vld(sys_arr_col4_vld[6]),
        .out1_data(sys_arr_col4_data[55:48]),
        .pe_doing(pe_doing[6][3]),
        .c1_vld(c1_vld[6][3]),
        .c1_data(c1_data[6][31:24])
    );
    
    pe u_pe_row6_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[4]),
        .in0_data(sys_arr_row6_data[39:32]),
        .in1_vld(sys_arr_col4_vld[6]),
        .in1_data(sys_arr_col4_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[4]),
        .out0_data(sys_arr_row7_data[39:32]),
        .out1_vld(sys_arr_col5_vld[6]),
        .out1_data(sys_arr_col5_data[55:48]),
        .pe_doing(pe_doing[6][4]),
        .c1_vld(c1_vld[6][4]),
        .c1_data(c1_data[6][39:32])
    );
    
    pe u_pe_row6_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[5]),
        .in0_data(sys_arr_row6_data[47:40]),
        .in1_vld(sys_arr_col5_vld[6]),
        .in1_data(sys_arr_col5_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[5]),
        .out0_data(sys_arr_row7_data[47:40]),
        .out1_vld(sys_arr_col6_vld[6]),
        .out1_data(sys_arr_col6_data[55:48]),
        .pe_doing(pe_doing[6][5]),
        .c1_vld(c1_vld[6][5]),
        .c1_data(c1_data[6][47:40])
    );
    
    pe u_pe_row6_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[6]),
        .in0_data(sys_arr_row6_data[55:48]),
        .in1_vld(sys_arr_col6_vld[6]),
        .in1_data(sys_arr_col6_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[6]),
        .out0_data(sys_arr_row7_data[55:48]),
        .out1_vld(sys_arr_col7_vld[6]),
        .out1_data(sys_arr_col7_data[55:48]),
        .pe_doing(pe_doing[6][6]),
        .c1_vld(c1_vld[6][6]),
        .c1_data(c1_data[6][55:48])
    );
    
    pe u_pe_row6_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[7]),
        .in0_data(sys_arr_row6_data[63:56]),
        .in1_vld(sys_arr_col7_vld[6]),
        .in1_data(sys_arr_col7_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[7]),
        .out0_data(sys_arr_row7_data[63:56]),
        .out1_vld(sys_arr_col8_vld[6]),
        .out1_data(sys_arr_col8_data[55:48]),
        .pe_doing(pe_doing[6][7]),
        .c1_vld(c1_vld[6][7]),
        .c1_data(c1_data[6][63:56])
    );
    
    pe u_pe_row6_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[8]),
        .in0_data(sys_arr_row6_data[71:64]),
        .in1_vld(sys_arr_col8_vld[6]),
        .in1_data(sys_arr_col8_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[8]),
        .out0_data(sys_arr_row7_data[71:64]),
        .out1_vld(sys_arr_col9_vld[6]),
        .out1_data(sys_arr_col9_data[55:48]),
        .pe_doing(pe_doing[6][8]),
        .c1_vld(c1_vld[6][8]),
        .c1_data(c1_data[6][71:64])
    );
    
    pe u_pe_row6_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[9]),
        .in0_data(sys_arr_row6_data[79:72]),
        .in1_vld(sys_arr_col9_vld[6]),
        .in1_data(sys_arr_col9_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[9]),
        .out0_data(sys_arr_row7_data[79:72]),
        .out1_vld(sys_arr_col10_vld[6]),
        .out1_data(sys_arr_col10_data[55:48]),
        .pe_doing(pe_doing[6][9]),
        .c1_vld(c1_vld[6][9]),
        .c1_data(c1_data[6][79:72])
    );
    
    pe u_pe_row6_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[10]),
        .in0_data(sys_arr_row6_data[87:80]),
        .in1_vld(sys_arr_col10_vld[6]),
        .in1_data(sys_arr_col10_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[10]),
        .out0_data(sys_arr_row7_data[87:80]),
        .out1_vld(sys_arr_col11_vld[6]),
        .out1_data(sys_arr_col11_data[55:48]),
        .pe_doing(pe_doing[6][10]),
        .c1_vld(c1_vld[6][10]),
        .c1_data(c1_data[6][87:80])
    );
    
    pe u_pe_row6_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[11]),
        .in0_data(sys_arr_row6_data[95:88]),
        .in1_vld(sys_arr_col11_vld[6]),
        .in1_data(sys_arr_col11_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[11]),
        .out0_data(sys_arr_row7_data[95:88]),
        .out1_vld(sys_arr_col12_vld[6]),
        .out1_data(sys_arr_col12_data[55:48]),
        .pe_doing(pe_doing[6][11]),
        .c1_vld(c1_vld[6][11]),
        .c1_data(c1_data[6][95:88])
    );
    
    pe u_pe_row6_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[12]),
        .in0_data(sys_arr_row6_data[103:96]),
        .in1_vld(sys_arr_col12_vld[6]),
        .in1_data(sys_arr_col12_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[12]),
        .out0_data(sys_arr_row7_data[103:96]),
        .out1_vld(sys_arr_col13_vld[6]),
        .out1_data(sys_arr_col13_data[55:48]),
        .pe_doing(pe_doing[6][12]),
        .c1_vld(c1_vld[6][12]),
        .c1_data(c1_data[6][103:96])
    );
    
    pe u_pe_row6_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[13]),
        .in0_data(sys_arr_row6_data[111:104]),
        .in1_vld(sys_arr_col13_vld[6]),
        .in1_data(sys_arr_col13_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[13]),
        .out0_data(sys_arr_row7_data[111:104]),
        .out1_vld(sys_arr_col14_vld[6]),
        .out1_data(sys_arr_col14_data[55:48]),
        .pe_doing(pe_doing[6][13]),
        .c1_vld(c1_vld[6][13]),
        .c1_data(c1_data[6][111:104])
    );
    
    pe u_pe_row6_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[14]),
        .in0_data(sys_arr_row6_data[119:112]),
        .in1_vld(sys_arr_col14_vld[6]),
        .in1_data(sys_arr_col14_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[14]),
        .out0_data(sys_arr_row7_data[119:112]),
        .out1_vld(sys_arr_col15_vld[6]),
        .out1_data(sys_arr_col15_data[55:48]),
        .pe_doing(pe_doing[6][14]),
        .c1_vld(c1_vld[6][14]),
        .c1_data(c1_data[6][119:112])
    );
    
    pe u_pe_row6_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row6_vld[15]),
        .in0_data(sys_arr_row6_data[127:120]),
        .in1_vld(sys_arr_col15_vld[6]),
        .in1_data(sys_arr_col15_data[55:48]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row7_vld[15]),
        .out0_data(sys_arr_row7_data[127:120]),
        .out1_vld(sys_arr_col16_vld[6]),
        .out1_data(sys_arr_col16_data[55:48]),
        .pe_doing(pe_doing[6][15]),
        .c1_vld(c1_vld[6][15]),
        .c1_data(c1_data[6][127:120])
    );
    
    pe u_pe_row7_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[0]),
        .in0_data(sys_arr_row7_data[7:0]),
        .in1_vld(sys_arr_col0_vld[7]),
        .in1_data(sys_arr_col0_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[0]),
        .out0_data(sys_arr_row8_data[7:0]),
        .out1_vld(sys_arr_col1_vld[7]),
        .out1_data(sys_arr_col1_data[63:56]),
        .pe_doing(pe_doing[7][0]),
        .c1_vld(c1_vld[7][0]),
        .c1_data(c1_data[7][7:0])
    );
    
    pe u_pe_row7_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[1]),
        .in0_data(sys_arr_row7_data[15:8]),
        .in1_vld(sys_arr_col1_vld[7]),
        .in1_data(sys_arr_col1_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[1]),
        .out0_data(sys_arr_row8_data[15:8]),
        .out1_vld(sys_arr_col2_vld[7]),
        .out1_data(sys_arr_col2_data[63:56]),
        .pe_doing(pe_doing[7][1]),
        .c1_vld(c1_vld[7][1]),
        .c1_data(c1_data[7][15:8])
    );
    
    pe u_pe_row7_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[2]),
        .in0_data(sys_arr_row7_data[23:16]),
        .in1_vld(sys_arr_col2_vld[7]),
        .in1_data(sys_arr_col2_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[2]),
        .out0_data(sys_arr_row8_data[23:16]),
        .out1_vld(sys_arr_col3_vld[7]),
        .out1_data(sys_arr_col3_data[63:56]),
        .pe_doing(pe_doing[7][2]),
        .c1_vld(c1_vld[7][2]),
        .c1_data(c1_data[7][23:16])
    );
    
    pe u_pe_row7_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[3]),
        .in0_data(sys_arr_row7_data[31:24]),
        .in1_vld(sys_arr_col3_vld[7]),
        .in1_data(sys_arr_col3_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[3]),
        .out0_data(sys_arr_row8_data[31:24]),
        .out1_vld(sys_arr_col4_vld[7]),
        .out1_data(sys_arr_col4_data[63:56]),
        .pe_doing(pe_doing[7][3]),
        .c1_vld(c1_vld[7][3]),
        .c1_data(c1_data[7][31:24])
    );
    
    pe u_pe_row7_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[4]),
        .in0_data(sys_arr_row7_data[39:32]),
        .in1_vld(sys_arr_col4_vld[7]),
        .in1_data(sys_arr_col4_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[4]),
        .out0_data(sys_arr_row8_data[39:32]),
        .out1_vld(sys_arr_col5_vld[7]),
        .out1_data(sys_arr_col5_data[63:56]),
        .pe_doing(pe_doing[7][4]),
        .c1_vld(c1_vld[7][4]),
        .c1_data(c1_data[7][39:32])
    );
    
    pe u_pe_row7_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[5]),
        .in0_data(sys_arr_row7_data[47:40]),
        .in1_vld(sys_arr_col5_vld[7]),
        .in1_data(sys_arr_col5_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[5]),
        .out0_data(sys_arr_row8_data[47:40]),
        .out1_vld(sys_arr_col6_vld[7]),
        .out1_data(sys_arr_col6_data[63:56]),
        .pe_doing(pe_doing[7][5]),
        .c1_vld(c1_vld[7][5]),
        .c1_data(c1_data[7][47:40])
    );
    
    pe u_pe_row7_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[6]),
        .in0_data(sys_arr_row7_data[55:48]),
        .in1_vld(sys_arr_col6_vld[7]),
        .in1_data(sys_arr_col6_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[6]),
        .out0_data(sys_arr_row8_data[55:48]),
        .out1_vld(sys_arr_col7_vld[7]),
        .out1_data(sys_arr_col7_data[63:56]),
        .pe_doing(pe_doing[7][6]),
        .c1_vld(c1_vld[7][6]),
        .c1_data(c1_data[7][55:48])
    );
    
    pe u_pe_row7_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[7]),
        .in0_data(sys_arr_row7_data[63:56]),
        .in1_vld(sys_arr_col7_vld[7]),
        .in1_data(sys_arr_col7_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[7]),
        .out0_data(sys_arr_row8_data[63:56]),
        .out1_vld(sys_arr_col8_vld[7]),
        .out1_data(sys_arr_col8_data[63:56]),
        .pe_doing(pe_doing[7][7]),
        .c1_vld(c1_vld[7][7]),
        .c1_data(c1_data[7][63:56])
    );
    
    pe u_pe_row7_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[8]),
        .in0_data(sys_arr_row7_data[71:64]),
        .in1_vld(sys_arr_col8_vld[7]),
        .in1_data(sys_arr_col8_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[8]),
        .out0_data(sys_arr_row8_data[71:64]),
        .out1_vld(sys_arr_col9_vld[7]),
        .out1_data(sys_arr_col9_data[63:56]),
        .pe_doing(pe_doing[7][8]),
        .c1_vld(c1_vld[7][8]),
        .c1_data(c1_data[7][71:64])
    );
    
    pe u_pe_row7_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[9]),
        .in0_data(sys_arr_row7_data[79:72]),
        .in1_vld(sys_arr_col9_vld[7]),
        .in1_data(sys_arr_col9_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[9]),
        .out0_data(sys_arr_row8_data[79:72]),
        .out1_vld(sys_arr_col10_vld[7]),
        .out1_data(sys_arr_col10_data[63:56]),
        .pe_doing(pe_doing[7][9]),
        .c1_vld(c1_vld[7][9]),
        .c1_data(c1_data[7][79:72])
    );
    
    pe u_pe_row7_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[10]),
        .in0_data(sys_arr_row7_data[87:80]),
        .in1_vld(sys_arr_col10_vld[7]),
        .in1_data(sys_arr_col10_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[10]),
        .out0_data(sys_arr_row8_data[87:80]),
        .out1_vld(sys_arr_col11_vld[7]),
        .out1_data(sys_arr_col11_data[63:56]),
        .pe_doing(pe_doing[7][10]),
        .c1_vld(c1_vld[7][10]),
        .c1_data(c1_data[7][87:80])
    );
    
    pe u_pe_row7_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[11]),
        .in0_data(sys_arr_row7_data[95:88]),
        .in1_vld(sys_arr_col11_vld[7]),
        .in1_data(sys_arr_col11_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[11]),
        .out0_data(sys_arr_row8_data[95:88]),
        .out1_vld(sys_arr_col12_vld[7]),
        .out1_data(sys_arr_col12_data[63:56]),
        .pe_doing(pe_doing[7][11]),
        .c1_vld(c1_vld[7][11]),
        .c1_data(c1_data[7][95:88])
    );
    
    pe u_pe_row7_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[12]),
        .in0_data(sys_arr_row7_data[103:96]),
        .in1_vld(sys_arr_col12_vld[7]),
        .in1_data(sys_arr_col12_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[12]),
        .out0_data(sys_arr_row8_data[103:96]),
        .out1_vld(sys_arr_col13_vld[7]),
        .out1_data(sys_arr_col13_data[63:56]),
        .pe_doing(pe_doing[7][12]),
        .c1_vld(c1_vld[7][12]),
        .c1_data(c1_data[7][103:96])
    );
    
    pe u_pe_row7_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[13]),
        .in0_data(sys_arr_row7_data[111:104]),
        .in1_vld(sys_arr_col13_vld[7]),
        .in1_data(sys_arr_col13_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[13]),
        .out0_data(sys_arr_row8_data[111:104]),
        .out1_vld(sys_arr_col14_vld[7]),
        .out1_data(sys_arr_col14_data[63:56]),
        .pe_doing(pe_doing[7][13]),
        .c1_vld(c1_vld[7][13]),
        .c1_data(c1_data[7][111:104])
    );
    
    pe u_pe_row7_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[14]),
        .in0_data(sys_arr_row7_data[119:112]),
        .in1_vld(sys_arr_col14_vld[7]),
        .in1_data(sys_arr_col14_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[14]),
        .out0_data(sys_arr_row8_data[119:112]),
        .out1_vld(sys_arr_col15_vld[7]),
        .out1_data(sys_arr_col15_data[63:56]),
        .pe_doing(pe_doing[7][14]),
        .c1_vld(c1_vld[7][14]),
        .c1_data(c1_data[7][119:112])
    );
    
    pe u_pe_row7_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row7_vld[15]),
        .in0_data(sys_arr_row7_data[127:120]),
        .in1_vld(sys_arr_col15_vld[7]),
        .in1_data(sys_arr_col15_data[63:56]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row8_vld[15]),
        .out0_data(sys_arr_row8_data[127:120]),
        .out1_vld(sys_arr_col16_vld[7]),
        .out1_data(sys_arr_col16_data[63:56]),
        .pe_doing(pe_doing[7][15]),
        .c1_vld(c1_vld[7][15]),
        .c1_data(c1_data[7][127:120])
    );
    
    pe u_pe_row8_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[0]),
        .in0_data(sys_arr_row8_data[7:0]),
        .in1_vld(sys_arr_col0_vld[8]),
        .in1_data(sys_arr_col0_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[0]),
        .out0_data(sys_arr_row9_data[7:0]),
        .out1_vld(sys_arr_col1_vld[8]),
        .out1_data(sys_arr_col1_data[71:64]),
        .pe_doing(pe_doing[8][0]),
        .c1_vld(c1_vld[8][0]),
        .c1_data(c1_data[8][7:0])
    );
    
    pe u_pe_row8_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[1]),
        .in0_data(sys_arr_row8_data[15:8]),
        .in1_vld(sys_arr_col1_vld[8]),
        .in1_data(sys_arr_col1_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[1]),
        .out0_data(sys_arr_row9_data[15:8]),
        .out1_vld(sys_arr_col2_vld[8]),
        .out1_data(sys_arr_col2_data[71:64]),
        .pe_doing(pe_doing[8][1]),
        .c1_vld(c1_vld[8][1]),
        .c1_data(c1_data[8][15:8])
    );
    
    pe u_pe_row8_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[2]),
        .in0_data(sys_arr_row8_data[23:16]),
        .in1_vld(sys_arr_col2_vld[8]),
        .in1_data(sys_arr_col2_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[2]),
        .out0_data(sys_arr_row9_data[23:16]),
        .out1_vld(sys_arr_col3_vld[8]),
        .out1_data(sys_arr_col3_data[71:64]),
        .pe_doing(pe_doing[8][2]),
        .c1_vld(c1_vld[8][2]),
        .c1_data(c1_data[8][23:16])
    );
    
    pe u_pe_row8_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[3]),
        .in0_data(sys_arr_row8_data[31:24]),
        .in1_vld(sys_arr_col3_vld[8]),
        .in1_data(sys_arr_col3_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[3]),
        .out0_data(sys_arr_row9_data[31:24]),
        .out1_vld(sys_arr_col4_vld[8]),
        .out1_data(sys_arr_col4_data[71:64]),
        .pe_doing(pe_doing[8][3]),
        .c1_vld(c1_vld[8][3]),
        .c1_data(c1_data[8][31:24])
    );
    
    pe u_pe_row8_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[4]),
        .in0_data(sys_arr_row8_data[39:32]),
        .in1_vld(sys_arr_col4_vld[8]),
        .in1_data(sys_arr_col4_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[4]),
        .out0_data(sys_arr_row9_data[39:32]),
        .out1_vld(sys_arr_col5_vld[8]),
        .out1_data(sys_arr_col5_data[71:64]),
        .pe_doing(pe_doing[8][4]),
        .c1_vld(c1_vld[8][4]),
        .c1_data(c1_data[8][39:32])
    );
    
    pe u_pe_row8_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[5]),
        .in0_data(sys_arr_row8_data[47:40]),
        .in1_vld(sys_arr_col5_vld[8]),
        .in1_data(sys_arr_col5_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[5]),
        .out0_data(sys_arr_row9_data[47:40]),
        .out1_vld(sys_arr_col6_vld[8]),
        .out1_data(sys_arr_col6_data[71:64]),
        .pe_doing(pe_doing[8][5]),
        .c1_vld(c1_vld[8][5]),
        .c1_data(c1_data[8][47:40])
    );
    
    pe u_pe_row8_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[6]),
        .in0_data(sys_arr_row8_data[55:48]),
        .in1_vld(sys_arr_col6_vld[8]),
        .in1_data(sys_arr_col6_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[6]),
        .out0_data(sys_arr_row9_data[55:48]),
        .out1_vld(sys_arr_col7_vld[8]),
        .out1_data(sys_arr_col7_data[71:64]),
        .pe_doing(pe_doing[8][6]),
        .c1_vld(c1_vld[8][6]),
        .c1_data(c1_data[8][55:48])
    );
    
    pe u_pe_row8_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[7]),
        .in0_data(sys_arr_row8_data[63:56]),
        .in1_vld(sys_arr_col7_vld[8]),
        .in1_data(sys_arr_col7_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[7]),
        .out0_data(sys_arr_row9_data[63:56]),
        .out1_vld(sys_arr_col8_vld[8]),
        .out1_data(sys_arr_col8_data[71:64]),
        .pe_doing(pe_doing[8][7]),
        .c1_vld(c1_vld[8][7]),
        .c1_data(c1_data[8][63:56])
    );
    
    pe u_pe_row8_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[8]),
        .in0_data(sys_arr_row8_data[71:64]),
        .in1_vld(sys_arr_col8_vld[8]),
        .in1_data(sys_arr_col8_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[8]),
        .out0_data(sys_arr_row9_data[71:64]),
        .out1_vld(sys_arr_col9_vld[8]),
        .out1_data(sys_arr_col9_data[71:64]),
        .pe_doing(pe_doing[8][8]),
        .c1_vld(c1_vld[8][8]),
        .c1_data(c1_data[8][71:64])
    );
    
    pe u_pe_row8_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[9]),
        .in0_data(sys_arr_row8_data[79:72]),
        .in1_vld(sys_arr_col9_vld[8]),
        .in1_data(sys_arr_col9_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[9]),
        .out0_data(sys_arr_row9_data[79:72]),
        .out1_vld(sys_arr_col10_vld[8]),
        .out1_data(sys_arr_col10_data[71:64]),
        .pe_doing(pe_doing[8][9]),
        .c1_vld(c1_vld[8][9]),
        .c1_data(c1_data[8][79:72])
    );
    
    pe u_pe_row8_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[10]),
        .in0_data(sys_arr_row8_data[87:80]),
        .in1_vld(sys_arr_col10_vld[8]),
        .in1_data(sys_arr_col10_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[10]),
        .out0_data(sys_arr_row9_data[87:80]),
        .out1_vld(sys_arr_col11_vld[8]),
        .out1_data(sys_arr_col11_data[71:64]),
        .pe_doing(pe_doing[8][10]),
        .c1_vld(c1_vld[8][10]),
        .c1_data(c1_data[8][87:80])
    );
    
    pe u_pe_row8_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[11]),
        .in0_data(sys_arr_row8_data[95:88]),
        .in1_vld(sys_arr_col11_vld[8]),
        .in1_data(sys_arr_col11_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[11]),
        .out0_data(sys_arr_row9_data[95:88]),
        .out1_vld(sys_arr_col12_vld[8]),
        .out1_data(sys_arr_col12_data[71:64]),
        .pe_doing(pe_doing[8][11]),
        .c1_vld(c1_vld[8][11]),
        .c1_data(c1_data[8][95:88])
    );
    
    pe u_pe_row8_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[12]),
        .in0_data(sys_arr_row8_data[103:96]),
        .in1_vld(sys_arr_col12_vld[8]),
        .in1_data(sys_arr_col12_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[12]),
        .out0_data(sys_arr_row9_data[103:96]),
        .out1_vld(sys_arr_col13_vld[8]),
        .out1_data(sys_arr_col13_data[71:64]),
        .pe_doing(pe_doing[8][12]),
        .c1_vld(c1_vld[8][12]),
        .c1_data(c1_data[8][103:96])
    );
    
    pe u_pe_row8_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[13]),
        .in0_data(sys_arr_row8_data[111:104]),
        .in1_vld(sys_arr_col13_vld[8]),
        .in1_data(sys_arr_col13_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[13]),
        .out0_data(sys_arr_row9_data[111:104]),
        .out1_vld(sys_arr_col14_vld[8]),
        .out1_data(sys_arr_col14_data[71:64]),
        .pe_doing(pe_doing[8][13]),
        .c1_vld(c1_vld[8][13]),
        .c1_data(c1_data[8][111:104])
    );
    
    pe u_pe_row8_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[14]),
        .in0_data(sys_arr_row8_data[119:112]),
        .in1_vld(sys_arr_col14_vld[8]),
        .in1_data(sys_arr_col14_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[14]),
        .out0_data(sys_arr_row9_data[119:112]),
        .out1_vld(sys_arr_col15_vld[8]),
        .out1_data(sys_arr_col15_data[71:64]),
        .pe_doing(pe_doing[8][14]),
        .c1_vld(c1_vld[8][14]),
        .c1_data(c1_data[8][119:112])
    );
    
    pe u_pe_row8_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row8_vld[15]),
        .in0_data(sys_arr_row8_data[127:120]),
        .in1_vld(sys_arr_col15_vld[8]),
        .in1_data(sys_arr_col15_data[71:64]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row9_vld[15]),
        .out0_data(sys_arr_row9_data[127:120]),
        .out1_vld(sys_arr_col16_vld[8]),
        .out1_data(sys_arr_col16_data[71:64]),
        .pe_doing(pe_doing[8][15]),
        .c1_vld(c1_vld[8][15]),
        .c1_data(c1_data[8][127:120])
    );
    
    pe u_pe_row9_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[0]),
        .in0_data(sys_arr_row9_data[7:0]),
        .in1_vld(sys_arr_col0_vld[9]),
        .in1_data(sys_arr_col0_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[0]),
        .out0_data(sys_arr_row10_data[7:0]),
        .out1_vld(sys_arr_col1_vld[9]),
        .out1_data(sys_arr_col1_data[79:72]),
        .pe_doing(pe_doing[9][0]),
        .c1_vld(c1_vld[9][0]),
        .c1_data(c1_data[9][7:0])
    );
    
    pe u_pe_row9_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[1]),
        .in0_data(sys_arr_row9_data[15:8]),
        .in1_vld(sys_arr_col1_vld[9]),
        .in1_data(sys_arr_col1_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[1]),
        .out0_data(sys_arr_row10_data[15:8]),
        .out1_vld(sys_arr_col2_vld[9]),
        .out1_data(sys_arr_col2_data[79:72]),
        .pe_doing(pe_doing[9][1]),
        .c1_vld(c1_vld[9][1]),
        .c1_data(c1_data[9][15:8])
    );
    
    pe u_pe_row9_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[2]),
        .in0_data(sys_arr_row9_data[23:16]),
        .in1_vld(sys_arr_col2_vld[9]),
        .in1_data(sys_arr_col2_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[2]),
        .out0_data(sys_arr_row10_data[23:16]),
        .out1_vld(sys_arr_col3_vld[9]),
        .out1_data(sys_arr_col3_data[79:72]),
        .pe_doing(pe_doing[9][2]),
        .c1_vld(c1_vld[9][2]),
        .c1_data(c1_data[9][23:16])
    );
    
    pe u_pe_row9_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[3]),
        .in0_data(sys_arr_row9_data[31:24]),
        .in1_vld(sys_arr_col3_vld[9]),
        .in1_data(sys_arr_col3_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[3]),
        .out0_data(sys_arr_row10_data[31:24]),
        .out1_vld(sys_arr_col4_vld[9]),
        .out1_data(sys_arr_col4_data[79:72]),
        .pe_doing(pe_doing[9][3]),
        .c1_vld(c1_vld[9][3]),
        .c1_data(c1_data[9][31:24])
    );
    
    pe u_pe_row9_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[4]),
        .in0_data(sys_arr_row9_data[39:32]),
        .in1_vld(sys_arr_col4_vld[9]),
        .in1_data(sys_arr_col4_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[4]),
        .out0_data(sys_arr_row10_data[39:32]),
        .out1_vld(sys_arr_col5_vld[9]),
        .out1_data(sys_arr_col5_data[79:72]),
        .pe_doing(pe_doing[9][4]),
        .c1_vld(c1_vld[9][4]),
        .c1_data(c1_data[9][39:32])
    );
    
    pe u_pe_row9_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[5]),
        .in0_data(sys_arr_row9_data[47:40]),
        .in1_vld(sys_arr_col5_vld[9]),
        .in1_data(sys_arr_col5_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[5]),
        .out0_data(sys_arr_row10_data[47:40]),
        .out1_vld(sys_arr_col6_vld[9]),
        .out1_data(sys_arr_col6_data[79:72]),
        .pe_doing(pe_doing[9][5]),
        .c1_vld(c1_vld[9][5]),
        .c1_data(c1_data[9][47:40])
    );
    
    pe u_pe_row9_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[6]),
        .in0_data(sys_arr_row9_data[55:48]),
        .in1_vld(sys_arr_col6_vld[9]),
        .in1_data(sys_arr_col6_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[6]),
        .out0_data(sys_arr_row10_data[55:48]),
        .out1_vld(sys_arr_col7_vld[9]),
        .out1_data(sys_arr_col7_data[79:72]),
        .pe_doing(pe_doing[9][6]),
        .c1_vld(c1_vld[9][6]),
        .c1_data(c1_data[9][55:48])
    );
    
    pe u_pe_row9_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[7]),
        .in0_data(sys_arr_row9_data[63:56]),
        .in1_vld(sys_arr_col7_vld[9]),
        .in1_data(sys_arr_col7_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[7]),
        .out0_data(sys_arr_row10_data[63:56]),
        .out1_vld(sys_arr_col8_vld[9]),
        .out1_data(sys_arr_col8_data[79:72]),
        .pe_doing(pe_doing[9][7]),
        .c1_vld(c1_vld[9][7]),
        .c1_data(c1_data[9][63:56])
    );
    
    pe u_pe_row9_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[8]),
        .in0_data(sys_arr_row9_data[71:64]),
        .in1_vld(sys_arr_col8_vld[9]),
        .in1_data(sys_arr_col8_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[8]),
        .out0_data(sys_arr_row10_data[71:64]),
        .out1_vld(sys_arr_col9_vld[9]),
        .out1_data(sys_arr_col9_data[79:72]),
        .pe_doing(pe_doing[9][8]),
        .c1_vld(c1_vld[9][8]),
        .c1_data(c1_data[9][71:64])
    );
    
    pe u_pe_row9_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[9]),
        .in0_data(sys_arr_row9_data[79:72]),
        .in1_vld(sys_arr_col9_vld[9]),
        .in1_data(sys_arr_col9_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[9]),
        .out0_data(sys_arr_row10_data[79:72]),
        .out1_vld(sys_arr_col10_vld[9]),
        .out1_data(sys_arr_col10_data[79:72]),
        .pe_doing(pe_doing[9][9]),
        .c1_vld(c1_vld[9][9]),
        .c1_data(c1_data[9][79:72])
    );
    
    pe u_pe_row9_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[10]),
        .in0_data(sys_arr_row9_data[87:80]),
        .in1_vld(sys_arr_col10_vld[9]),
        .in1_data(sys_arr_col10_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[10]),
        .out0_data(sys_arr_row10_data[87:80]),
        .out1_vld(sys_arr_col11_vld[9]),
        .out1_data(sys_arr_col11_data[79:72]),
        .pe_doing(pe_doing[9][10]),
        .c1_vld(c1_vld[9][10]),
        .c1_data(c1_data[9][87:80])
    );
    
    pe u_pe_row9_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[11]),
        .in0_data(sys_arr_row9_data[95:88]),
        .in1_vld(sys_arr_col11_vld[9]),
        .in1_data(sys_arr_col11_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[11]),
        .out0_data(sys_arr_row10_data[95:88]),
        .out1_vld(sys_arr_col12_vld[9]),
        .out1_data(sys_arr_col12_data[79:72]),
        .pe_doing(pe_doing[9][11]),
        .c1_vld(c1_vld[9][11]),
        .c1_data(c1_data[9][95:88])
    );
    
    pe u_pe_row9_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[12]),
        .in0_data(sys_arr_row9_data[103:96]),
        .in1_vld(sys_arr_col12_vld[9]),
        .in1_data(sys_arr_col12_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[12]),
        .out0_data(sys_arr_row10_data[103:96]),
        .out1_vld(sys_arr_col13_vld[9]),
        .out1_data(sys_arr_col13_data[79:72]),
        .pe_doing(pe_doing[9][12]),
        .c1_vld(c1_vld[9][12]),
        .c1_data(c1_data[9][103:96])
    );
    
    pe u_pe_row9_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[13]),
        .in0_data(sys_arr_row9_data[111:104]),
        .in1_vld(sys_arr_col13_vld[9]),
        .in1_data(sys_arr_col13_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[13]),
        .out0_data(sys_arr_row10_data[111:104]),
        .out1_vld(sys_arr_col14_vld[9]),
        .out1_data(sys_arr_col14_data[79:72]),
        .pe_doing(pe_doing[9][13]),
        .c1_vld(c1_vld[9][13]),
        .c1_data(c1_data[9][111:104])
    );
    
    pe u_pe_row9_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[14]),
        .in0_data(sys_arr_row9_data[119:112]),
        .in1_vld(sys_arr_col14_vld[9]),
        .in1_data(sys_arr_col14_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[14]),
        .out0_data(sys_arr_row10_data[119:112]),
        .out1_vld(sys_arr_col15_vld[9]),
        .out1_data(sys_arr_col15_data[79:72]),
        .pe_doing(pe_doing[9][14]),
        .c1_vld(c1_vld[9][14]),
        .c1_data(c1_data[9][119:112])
    );
    
    pe u_pe_row9_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row9_vld[15]),
        .in0_data(sys_arr_row9_data[127:120]),
        .in1_vld(sys_arr_col15_vld[9]),
        .in1_data(sys_arr_col15_data[79:72]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row10_vld[15]),
        .out0_data(sys_arr_row10_data[127:120]),
        .out1_vld(sys_arr_col16_vld[9]),
        .out1_data(sys_arr_col16_data[79:72]),
        .pe_doing(pe_doing[9][15]),
        .c1_vld(c1_vld[9][15]),
        .c1_data(c1_data[9][127:120])
    );
    
    pe u_pe_row10_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[0]),
        .in0_data(sys_arr_row10_data[7:0]),
        .in1_vld(sys_arr_col0_vld[10]),
        .in1_data(sys_arr_col0_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[0]),
        .out0_data(sys_arr_row11_data[7:0]),
        .out1_vld(sys_arr_col1_vld[10]),
        .out1_data(sys_arr_col1_data[87:80]),
        .pe_doing(pe_doing[10][0]),
        .c1_vld(c1_vld[10][0]),
        .c1_data(c1_data[10][7:0])
    );
    
    pe u_pe_row10_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[1]),
        .in0_data(sys_arr_row10_data[15:8]),
        .in1_vld(sys_arr_col1_vld[10]),
        .in1_data(sys_arr_col1_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[1]),
        .out0_data(sys_arr_row11_data[15:8]),
        .out1_vld(sys_arr_col2_vld[10]),
        .out1_data(sys_arr_col2_data[87:80]),
        .pe_doing(pe_doing[10][1]),
        .c1_vld(c1_vld[10][1]),
        .c1_data(c1_data[10][15:8])
    );
    
    pe u_pe_row10_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[2]),
        .in0_data(sys_arr_row10_data[23:16]),
        .in1_vld(sys_arr_col2_vld[10]),
        .in1_data(sys_arr_col2_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[2]),
        .out0_data(sys_arr_row11_data[23:16]),
        .out1_vld(sys_arr_col3_vld[10]),
        .out1_data(sys_arr_col3_data[87:80]),
        .pe_doing(pe_doing[10][2]),
        .c1_vld(c1_vld[10][2]),
        .c1_data(c1_data[10][23:16])
    );
    
    pe u_pe_row10_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[3]),
        .in0_data(sys_arr_row10_data[31:24]),
        .in1_vld(sys_arr_col3_vld[10]),
        .in1_data(sys_arr_col3_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[3]),
        .out0_data(sys_arr_row11_data[31:24]),
        .out1_vld(sys_arr_col4_vld[10]),
        .out1_data(sys_arr_col4_data[87:80]),
        .pe_doing(pe_doing[10][3]),
        .c1_vld(c1_vld[10][3]),
        .c1_data(c1_data[10][31:24])
    );
    
    pe u_pe_row10_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[4]),
        .in0_data(sys_arr_row10_data[39:32]),
        .in1_vld(sys_arr_col4_vld[10]),
        .in1_data(sys_arr_col4_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[4]),
        .out0_data(sys_arr_row11_data[39:32]),
        .out1_vld(sys_arr_col5_vld[10]),
        .out1_data(sys_arr_col5_data[87:80]),
        .pe_doing(pe_doing[10][4]),
        .c1_vld(c1_vld[10][4]),
        .c1_data(c1_data[10][39:32])
    );
    
    pe u_pe_row10_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[5]),
        .in0_data(sys_arr_row10_data[47:40]),
        .in1_vld(sys_arr_col5_vld[10]),
        .in1_data(sys_arr_col5_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[5]),
        .out0_data(sys_arr_row11_data[47:40]),
        .out1_vld(sys_arr_col6_vld[10]),
        .out1_data(sys_arr_col6_data[87:80]),
        .pe_doing(pe_doing[10][5]),
        .c1_vld(c1_vld[10][5]),
        .c1_data(c1_data[10][47:40])
    );
    
    pe u_pe_row10_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[6]),
        .in0_data(sys_arr_row10_data[55:48]),
        .in1_vld(sys_arr_col6_vld[10]),
        .in1_data(sys_arr_col6_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[6]),
        .out0_data(sys_arr_row11_data[55:48]),
        .out1_vld(sys_arr_col7_vld[10]),
        .out1_data(sys_arr_col7_data[87:80]),
        .pe_doing(pe_doing[10][6]),
        .c1_vld(c1_vld[10][6]),
        .c1_data(c1_data[10][55:48])
    );
    
    pe u_pe_row10_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[7]),
        .in0_data(sys_arr_row10_data[63:56]),
        .in1_vld(sys_arr_col7_vld[10]),
        .in1_data(sys_arr_col7_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[7]),
        .out0_data(sys_arr_row11_data[63:56]),
        .out1_vld(sys_arr_col8_vld[10]),
        .out1_data(sys_arr_col8_data[87:80]),
        .pe_doing(pe_doing[10][7]),
        .c1_vld(c1_vld[10][7]),
        .c1_data(c1_data[10][63:56])
    );
    
    pe u_pe_row10_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[8]),
        .in0_data(sys_arr_row10_data[71:64]),
        .in1_vld(sys_arr_col8_vld[10]),
        .in1_data(sys_arr_col8_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[8]),
        .out0_data(sys_arr_row11_data[71:64]),
        .out1_vld(sys_arr_col9_vld[10]),
        .out1_data(sys_arr_col9_data[87:80]),
        .pe_doing(pe_doing[10][8]),
        .c1_vld(c1_vld[10][8]),
        .c1_data(c1_data[10][71:64])
    );
    
    pe u_pe_row10_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[9]),
        .in0_data(sys_arr_row10_data[79:72]),
        .in1_vld(sys_arr_col9_vld[10]),
        .in1_data(sys_arr_col9_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[9]),
        .out0_data(sys_arr_row11_data[79:72]),
        .out1_vld(sys_arr_col10_vld[10]),
        .out1_data(sys_arr_col10_data[87:80]),
        .pe_doing(pe_doing[10][9]),
        .c1_vld(c1_vld[10][9]),
        .c1_data(c1_data[10][79:72])
    );
    
    pe u_pe_row10_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[10]),
        .in0_data(sys_arr_row10_data[87:80]),
        .in1_vld(sys_arr_col10_vld[10]),
        .in1_data(sys_arr_col10_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[10]),
        .out0_data(sys_arr_row11_data[87:80]),
        .out1_vld(sys_arr_col11_vld[10]),
        .out1_data(sys_arr_col11_data[87:80]),
        .pe_doing(pe_doing[10][10]),
        .c1_vld(c1_vld[10][10]),
        .c1_data(c1_data[10][87:80])
    );
    
    pe u_pe_row10_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[11]),
        .in0_data(sys_arr_row10_data[95:88]),
        .in1_vld(sys_arr_col11_vld[10]),
        .in1_data(sys_arr_col11_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[11]),
        .out0_data(sys_arr_row11_data[95:88]),
        .out1_vld(sys_arr_col12_vld[10]),
        .out1_data(sys_arr_col12_data[87:80]),
        .pe_doing(pe_doing[10][11]),
        .c1_vld(c1_vld[10][11]),
        .c1_data(c1_data[10][95:88])
    );
    
    pe u_pe_row10_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[12]),
        .in0_data(sys_arr_row10_data[103:96]),
        .in1_vld(sys_arr_col12_vld[10]),
        .in1_data(sys_arr_col12_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[12]),
        .out0_data(sys_arr_row11_data[103:96]),
        .out1_vld(sys_arr_col13_vld[10]),
        .out1_data(sys_arr_col13_data[87:80]),
        .pe_doing(pe_doing[10][12]),
        .c1_vld(c1_vld[10][12]),
        .c1_data(c1_data[10][103:96])
    );
    
    pe u_pe_row10_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[13]),
        .in0_data(sys_arr_row10_data[111:104]),
        .in1_vld(sys_arr_col13_vld[10]),
        .in1_data(sys_arr_col13_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[13]),
        .out0_data(sys_arr_row11_data[111:104]),
        .out1_vld(sys_arr_col14_vld[10]),
        .out1_data(sys_arr_col14_data[87:80]),
        .pe_doing(pe_doing[10][13]),
        .c1_vld(c1_vld[10][13]),
        .c1_data(c1_data[10][111:104])
    );
    
    pe u_pe_row10_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[14]),
        .in0_data(sys_arr_row10_data[119:112]),
        .in1_vld(sys_arr_col14_vld[10]),
        .in1_data(sys_arr_col14_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[14]),
        .out0_data(sys_arr_row11_data[119:112]),
        .out1_vld(sys_arr_col15_vld[10]),
        .out1_data(sys_arr_col15_data[87:80]),
        .pe_doing(pe_doing[10][14]),
        .c1_vld(c1_vld[10][14]),
        .c1_data(c1_data[10][119:112])
    );
    
    pe u_pe_row10_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row10_vld[15]),
        .in0_data(sys_arr_row10_data[127:120]),
        .in1_vld(sys_arr_col15_vld[10]),
        .in1_data(sys_arr_col15_data[87:80]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row11_vld[15]),
        .out0_data(sys_arr_row11_data[127:120]),
        .out1_vld(sys_arr_col16_vld[10]),
        .out1_data(sys_arr_col16_data[87:80]),
        .pe_doing(pe_doing[10][15]),
        .c1_vld(c1_vld[10][15]),
        .c1_data(c1_data[10][127:120])
    );
    
    pe u_pe_row11_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[0]),
        .in0_data(sys_arr_row11_data[7:0]),
        .in1_vld(sys_arr_col0_vld[11]),
        .in1_data(sys_arr_col0_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[0]),
        .out0_data(sys_arr_row12_data[7:0]),
        .out1_vld(sys_arr_col1_vld[11]),
        .out1_data(sys_arr_col1_data[95:88]),
        .pe_doing(pe_doing[11][0]),
        .c1_vld(c1_vld[11][0]),
        .c1_data(c1_data[11][7:0])
    );
    
    pe u_pe_row11_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[1]),
        .in0_data(sys_arr_row11_data[15:8]),
        .in1_vld(sys_arr_col1_vld[11]),
        .in1_data(sys_arr_col1_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[1]),
        .out0_data(sys_arr_row12_data[15:8]),
        .out1_vld(sys_arr_col2_vld[11]),
        .out1_data(sys_arr_col2_data[95:88]),
        .pe_doing(pe_doing[11][1]),
        .c1_vld(c1_vld[11][1]),
        .c1_data(c1_data[11][15:8])
    );
    
    pe u_pe_row11_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[2]),
        .in0_data(sys_arr_row11_data[23:16]),
        .in1_vld(sys_arr_col2_vld[11]),
        .in1_data(sys_arr_col2_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[2]),
        .out0_data(sys_arr_row12_data[23:16]),
        .out1_vld(sys_arr_col3_vld[11]),
        .out1_data(sys_arr_col3_data[95:88]),
        .pe_doing(pe_doing[11][2]),
        .c1_vld(c1_vld[11][2]),
        .c1_data(c1_data[11][23:16])
    );
    
    pe u_pe_row11_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[3]),
        .in0_data(sys_arr_row11_data[31:24]),
        .in1_vld(sys_arr_col3_vld[11]),
        .in1_data(sys_arr_col3_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[3]),
        .out0_data(sys_arr_row12_data[31:24]),
        .out1_vld(sys_arr_col4_vld[11]),
        .out1_data(sys_arr_col4_data[95:88]),
        .pe_doing(pe_doing[11][3]),
        .c1_vld(c1_vld[11][3]),
        .c1_data(c1_data[11][31:24])
    );
    
    pe u_pe_row11_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[4]),
        .in0_data(sys_arr_row11_data[39:32]),
        .in1_vld(sys_arr_col4_vld[11]),
        .in1_data(sys_arr_col4_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[4]),
        .out0_data(sys_arr_row12_data[39:32]),
        .out1_vld(sys_arr_col5_vld[11]),
        .out1_data(sys_arr_col5_data[95:88]),
        .pe_doing(pe_doing[11][4]),
        .c1_vld(c1_vld[11][4]),
        .c1_data(c1_data[11][39:32])
    );
    
    pe u_pe_row11_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[5]),
        .in0_data(sys_arr_row11_data[47:40]),
        .in1_vld(sys_arr_col5_vld[11]),
        .in1_data(sys_arr_col5_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[5]),
        .out0_data(sys_arr_row12_data[47:40]),
        .out1_vld(sys_arr_col6_vld[11]),
        .out1_data(sys_arr_col6_data[95:88]),
        .pe_doing(pe_doing[11][5]),
        .c1_vld(c1_vld[11][5]),
        .c1_data(c1_data[11][47:40])
    );
    
    pe u_pe_row11_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[6]),
        .in0_data(sys_arr_row11_data[55:48]),
        .in1_vld(sys_arr_col6_vld[11]),
        .in1_data(sys_arr_col6_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[6]),
        .out0_data(sys_arr_row12_data[55:48]),
        .out1_vld(sys_arr_col7_vld[11]),
        .out1_data(sys_arr_col7_data[95:88]),
        .pe_doing(pe_doing[11][6]),
        .c1_vld(c1_vld[11][6]),
        .c1_data(c1_data[11][55:48])
    );
    
    pe u_pe_row11_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[7]),
        .in0_data(sys_arr_row11_data[63:56]),
        .in1_vld(sys_arr_col7_vld[11]),
        .in1_data(sys_arr_col7_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[7]),
        .out0_data(sys_arr_row12_data[63:56]),
        .out1_vld(sys_arr_col8_vld[11]),
        .out1_data(sys_arr_col8_data[95:88]),
        .pe_doing(pe_doing[11][7]),
        .c1_vld(c1_vld[11][7]),
        .c1_data(c1_data[11][63:56])
    );
    
    pe u_pe_row11_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[8]),
        .in0_data(sys_arr_row11_data[71:64]),
        .in1_vld(sys_arr_col8_vld[11]),
        .in1_data(sys_arr_col8_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[8]),
        .out0_data(sys_arr_row12_data[71:64]),
        .out1_vld(sys_arr_col9_vld[11]),
        .out1_data(sys_arr_col9_data[95:88]),
        .pe_doing(pe_doing[11][8]),
        .c1_vld(c1_vld[11][8]),
        .c1_data(c1_data[11][71:64])
    );
    
    pe u_pe_row11_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[9]),
        .in0_data(sys_arr_row11_data[79:72]),
        .in1_vld(sys_arr_col9_vld[11]),
        .in1_data(sys_arr_col9_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[9]),
        .out0_data(sys_arr_row12_data[79:72]),
        .out1_vld(sys_arr_col10_vld[11]),
        .out1_data(sys_arr_col10_data[95:88]),
        .pe_doing(pe_doing[11][9]),
        .c1_vld(c1_vld[11][9]),
        .c1_data(c1_data[11][79:72])
    );
    
    pe u_pe_row11_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[10]),
        .in0_data(sys_arr_row11_data[87:80]),
        .in1_vld(sys_arr_col10_vld[11]),
        .in1_data(sys_arr_col10_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[10]),
        .out0_data(sys_arr_row12_data[87:80]),
        .out1_vld(sys_arr_col11_vld[11]),
        .out1_data(sys_arr_col11_data[95:88]),
        .pe_doing(pe_doing[11][10]),
        .c1_vld(c1_vld[11][10]),
        .c1_data(c1_data[11][87:80])
    );
    
    pe u_pe_row11_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[11]),
        .in0_data(sys_arr_row11_data[95:88]),
        .in1_vld(sys_arr_col11_vld[11]),
        .in1_data(sys_arr_col11_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[11]),
        .out0_data(sys_arr_row12_data[95:88]),
        .out1_vld(sys_arr_col12_vld[11]),
        .out1_data(sys_arr_col12_data[95:88]),
        .pe_doing(pe_doing[11][11]),
        .c1_vld(c1_vld[11][11]),
        .c1_data(c1_data[11][95:88])
    );
    
    pe u_pe_row11_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[12]),
        .in0_data(sys_arr_row11_data[103:96]),
        .in1_vld(sys_arr_col12_vld[11]),
        .in1_data(sys_arr_col12_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[12]),
        .out0_data(sys_arr_row12_data[103:96]),
        .out1_vld(sys_arr_col13_vld[11]),
        .out1_data(sys_arr_col13_data[95:88]),
        .pe_doing(pe_doing[11][12]),
        .c1_vld(c1_vld[11][12]),
        .c1_data(c1_data[11][103:96])
    );
    
    pe u_pe_row11_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[13]),
        .in0_data(sys_arr_row11_data[111:104]),
        .in1_vld(sys_arr_col13_vld[11]),
        .in1_data(sys_arr_col13_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[13]),
        .out0_data(sys_arr_row12_data[111:104]),
        .out1_vld(sys_arr_col14_vld[11]),
        .out1_data(sys_arr_col14_data[95:88]),
        .pe_doing(pe_doing[11][13]),
        .c1_vld(c1_vld[11][13]),
        .c1_data(c1_data[11][111:104])
    );
    
    pe u_pe_row11_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[14]),
        .in0_data(sys_arr_row11_data[119:112]),
        .in1_vld(sys_arr_col14_vld[11]),
        .in1_data(sys_arr_col14_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[14]),
        .out0_data(sys_arr_row12_data[119:112]),
        .out1_vld(sys_arr_col15_vld[11]),
        .out1_data(sys_arr_col15_data[95:88]),
        .pe_doing(pe_doing[11][14]),
        .c1_vld(c1_vld[11][14]),
        .c1_data(c1_data[11][119:112])
    );
    
    pe u_pe_row11_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row11_vld[15]),
        .in0_data(sys_arr_row11_data[127:120]),
        .in1_vld(sys_arr_col15_vld[11]),
        .in1_data(sys_arr_col15_data[95:88]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row12_vld[15]),
        .out0_data(sys_arr_row12_data[127:120]),
        .out1_vld(sys_arr_col16_vld[11]),
        .out1_data(sys_arr_col16_data[95:88]),
        .pe_doing(pe_doing[11][15]),
        .c1_vld(c1_vld[11][15]),
        .c1_data(c1_data[11][127:120])
    );
    
    pe u_pe_row12_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[0]),
        .in0_data(sys_arr_row12_data[7:0]),
        .in1_vld(sys_arr_col0_vld[12]),
        .in1_data(sys_arr_col0_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[0]),
        .out0_data(sys_arr_row13_data[7:0]),
        .out1_vld(sys_arr_col1_vld[12]),
        .out1_data(sys_arr_col1_data[103:96]),
        .pe_doing(pe_doing[12][0]),
        .c1_vld(c1_vld[12][0]),
        .c1_data(c1_data[12][7:0])
    );
    
    pe u_pe_row12_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[1]),
        .in0_data(sys_arr_row12_data[15:8]),
        .in1_vld(sys_arr_col1_vld[12]),
        .in1_data(sys_arr_col1_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[1]),
        .out0_data(sys_arr_row13_data[15:8]),
        .out1_vld(sys_arr_col2_vld[12]),
        .out1_data(sys_arr_col2_data[103:96]),
        .pe_doing(pe_doing[12][1]),
        .c1_vld(c1_vld[12][1]),
        .c1_data(c1_data[12][15:8])
    );
    
    pe u_pe_row12_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[2]),
        .in0_data(sys_arr_row12_data[23:16]),
        .in1_vld(sys_arr_col2_vld[12]),
        .in1_data(sys_arr_col2_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[2]),
        .out0_data(sys_arr_row13_data[23:16]),
        .out1_vld(sys_arr_col3_vld[12]),
        .out1_data(sys_arr_col3_data[103:96]),
        .pe_doing(pe_doing[12][2]),
        .c1_vld(c1_vld[12][2]),
        .c1_data(c1_data[12][23:16])
    );
    
    pe u_pe_row12_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[3]),
        .in0_data(sys_arr_row12_data[31:24]),
        .in1_vld(sys_arr_col3_vld[12]),
        .in1_data(sys_arr_col3_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[3]),
        .out0_data(sys_arr_row13_data[31:24]),
        .out1_vld(sys_arr_col4_vld[12]),
        .out1_data(sys_arr_col4_data[103:96]),
        .pe_doing(pe_doing[12][3]),
        .c1_vld(c1_vld[12][3]),
        .c1_data(c1_data[12][31:24])
    );
    
    pe u_pe_row12_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[4]),
        .in0_data(sys_arr_row12_data[39:32]),
        .in1_vld(sys_arr_col4_vld[12]),
        .in1_data(sys_arr_col4_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[4]),
        .out0_data(sys_arr_row13_data[39:32]),
        .out1_vld(sys_arr_col5_vld[12]),
        .out1_data(sys_arr_col5_data[103:96]),
        .pe_doing(pe_doing[12][4]),
        .c1_vld(c1_vld[12][4]),
        .c1_data(c1_data[12][39:32])
    );
    
    pe u_pe_row12_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[5]),
        .in0_data(sys_arr_row12_data[47:40]),
        .in1_vld(sys_arr_col5_vld[12]),
        .in1_data(sys_arr_col5_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[5]),
        .out0_data(sys_arr_row13_data[47:40]),
        .out1_vld(sys_arr_col6_vld[12]),
        .out1_data(sys_arr_col6_data[103:96]),
        .pe_doing(pe_doing[12][5]),
        .c1_vld(c1_vld[12][5]),
        .c1_data(c1_data[12][47:40])
    );
    
    pe u_pe_row12_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[6]),
        .in0_data(sys_arr_row12_data[55:48]),
        .in1_vld(sys_arr_col6_vld[12]),
        .in1_data(sys_arr_col6_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[6]),
        .out0_data(sys_arr_row13_data[55:48]),
        .out1_vld(sys_arr_col7_vld[12]),
        .out1_data(sys_arr_col7_data[103:96]),
        .pe_doing(pe_doing[12][6]),
        .c1_vld(c1_vld[12][6]),
        .c1_data(c1_data[12][55:48])
    );
    
    pe u_pe_row12_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[7]),
        .in0_data(sys_arr_row12_data[63:56]),
        .in1_vld(sys_arr_col7_vld[12]),
        .in1_data(sys_arr_col7_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[7]),
        .out0_data(sys_arr_row13_data[63:56]),
        .out1_vld(sys_arr_col8_vld[12]),
        .out1_data(sys_arr_col8_data[103:96]),
        .pe_doing(pe_doing[12][7]),
        .c1_vld(c1_vld[12][7]),
        .c1_data(c1_data[12][63:56])
    );
    
    pe u_pe_row12_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[8]),
        .in0_data(sys_arr_row12_data[71:64]),
        .in1_vld(sys_arr_col8_vld[12]),
        .in1_data(sys_arr_col8_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[8]),
        .out0_data(sys_arr_row13_data[71:64]),
        .out1_vld(sys_arr_col9_vld[12]),
        .out1_data(sys_arr_col9_data[103:96]),
        .pe_doing(pe_doing[12][8]),
        .c1_vld(c1_vld[12][8]),
        .c1_data(c1_data[12][71:64])
    );
    
    pe u_pe_row12_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[9]),
        .in0_data(sys_arr_row12_data[79:72]),
        .in1_vld(sys_arr_col9_vld[12]),
        .in1_data(sys_arr_col9_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[9]),
        .out0_data(sys_arr_row13_data[79:72]),
        .out1_vld(sys_arr_col10_vld[12]),
        .out1_data(sys_arr_col10_data[103:96]),
        .pe_doing(pe_doing[12][9]),
        .c1_vld(c1_vld[12][9]),
        .c1_data(c1_data[12][79:72])
    );
    
    pe u_pe_row12_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[10]),
        .in0_data(sys_arr_row12_data[87:80]),
        .in1_vld(sys_arr_col10_vld[12]),
        .in1_data(sys_arr_col10_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[10]),
        .out0_data(sys_arr_row13_data[87:80]),
        .out1_vld(sys_arr_col11_vld[12]),
        .out1_data(sys_arr_col11_data[103:96]),
        .pe_doing(pe_doing[12][10]),
        .c1_vld(c1_vld[12][10]),
        .c1_data(c1_data[12][87:80])
    );
    
    pe u_pe_row12_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[11]),
        .in0_data(sys_arr_row12_data[95:88]),
        .in1_vld(sys_arr_col11_vld[12]),
        .in1_data(sys_arr_col11_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[11]),
        .out0_data(sys_arr_row13_data[95:88]),
        .out1_vld(sys_arr_col12_vld[12]),
        .out1_data(sys_arr_col12_data[103:96]),
        .pe_doing(pe_doing[12][11]),
        .c1_vld(c1_vld[12][11]),
        .c1_data(c1_data[12][95:88])
    );
    
    pe u_pe_row12_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[12]),
        .in0_data(sys_arr_row12_data[103:96]),
        .in1_vld(sys_arr_col12_vld[12]),
        .in1_data(sys_arr_col12_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[12]),
        .out0_data(sys_arr_row13_data[103:96]),
        .out1_vld(sys_arr_col13_vld[12]),
        .out1_data(sys_arr_col13_data[103:96]),
        .pe_doing(pe_doing[12][12]),
        .c1_vld(c1_vld[12][12]),
        .c1_data(c1_data[12][103:96])
    );
    
    pe u_pe_row12_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[13]),
        .in0_data(sys_arr_row12_data[111:104]),
        .in1_vld(sys_arr_col13_vld[12]),
        .in1_data(sys_arr_col13_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[13]),
        .out0_data(sys_arr_row13_data[111:104]),
        .out1_vld(sys_arr_col14_vld[12]),
        .out1_data(sys_arr_col14_data[103:96]),
        .pe_doing(pe_doing[12][13]),
        .c1_vld(c1_vld[12][13]),
        .c1_data(c1_data[12][111:104])
    );
    
    pe u_pe_row12_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[14]),
        .in0_data(sys_arr_row12_data[119:112]),
        .in1_vld(sys_arr_col14_vld[12]),
        .in1_data(sys_arr_col14_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[14]),
        .out0_data(sys_arr_row13_data[119:112]),
        .out1_vld(sys_arr_col15_vld[12]),
        .out1_data(sys_arr_col15_data[103:96]),
        .pe_doing(pe_doing[12][14]),
        .c1_vld(c1_vld[12][14]),
        .c1_data(c1_data[12][119:112])
    );
    
    pe u_pe_row12_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row12_vld[15]),
        .in0_data(sys_arr_row12_data[127:120]),
        .in1_vld(sys_arr_col15_vld[12]),
        .in1_data(sys_arr_col15_data[103:96]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row13_vld[15]),
        .out0_data(sys_arr_row13_data[127:120]),
        .out1_vld(sys_arr_col16_vld[12]),
        .out1_data(sys_arr_col16_data[103:96]),
        .pe_doing(pe_doing[12][15]),
        .c1_vld(c1_vld[12][15]),
        .c1_data(c1_data[12][127:120])
    );
    
    pe u_pe_row13_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[0]),
        .in0_data(sys_arr_row13_data[7:0]),
        .in1_vld(sys_arr_col0_vld[13]),
        .in1_data(sys_arr_col0_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[0]),
        .out0_data(sys_arr_row14_data[7:0]),
        .out1_vld(sys_arr_col1_vld[13]),
        .out1_data(sys_arr_col1_data[111:104]),
        .pe_doing(pe_doing[13][0]),
        .c1_vld(c1_vld[13][0]),
        .c1_data(c1_data[13][7:0])
    );
    
    pe u_pe_row13_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[1]),
        .in0_data(sys_arr_row13_data[15:8]),
        .in1_vld(sys_arr_col1_vld[13]),
        .in1_data(sys_arr_col1_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[1]),
        .out0_data(sys_arr_row14_data[15:8]),
        .out1_vld(sys_arr_col2_vld[13]),
        .out1_data(sys_arr_col2_data[111:104]),
        .pe_doing(pe_doing[13][1]),
        .c1_vld(c1_vld[13][1]),
        .c1_data(c1_data[13][15:8])
    );
    
    pe u_pe_row13_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[2]),
        .in0_data(sys_arr_row13_data[23:16]),
        .in1_vld(sys_arr_col2_vld[13]),
        .in1_data(sys_arr_col2_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[2]),
        .out0_data(sys_arr_row14_data[23:16]),
        .out1_vld(sys_arr_col3_vld[13]),
        .out1_data(sys_arr_col3_data[111:104]),
        .pe_doing(pe_doing[13][2]),
        .c1_vld(c1_vld[13][2]),
        .c1_data(c1_data[13][23:16])
    );
    
    pe u_pe_row13_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[3]),
        .in0_data(sys_arr_row13_data[31:24]),
        .in1_vld(sys_arr_col3_vld[13]),
        .in1_data(sys_arr_col3_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[3]),
        .out0_data(sys_arr_row14_data[31:24]),
        .out1_vld(sys_arr_col4_vld[13]),
        .out1_data(sys_arr_col4_data[111:104]),
        .pe_doing(pe_doing[13][3]),
        .c1_vld(c1_vld[13][3]),
        .c1_data(c1_data[13][31:24])
    );
    
    pe u_pe_row13_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[4]),
        .in0_data(sys_arr_row13_data[39:32]),
        .in1_vld(sys_arr_col4_vld[13]),
        .in1_data(sys_arr_col4_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[4]),
        .out0_data(sys_arr_row14_data[39:32]),
        .out1_vld(sys_arr_col5_vld[13]),
        .out1_data(sys_arr_col5_data[111:104]),
        .pe_doing(pe_doing[13][4]),
        .c1_vld(c1_vld[13][4]),
        .c1_data(c1_data[13][39:32])
    );
    
    pe u_pe_row13_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[5]),
        .in0_data(sys_arr_row13_data[47:40]),
        .in1_vld(sys_arr_col5_vld[13]),
        .in1_data(sys_arr_col5_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[5]),
        .out0_data(sys_arr_row14_data[47:40]),
        .out1_vld(sys_arr_col6_vld[13]),
        .out1_data(sys_arr_col6_data[111:104]),
        .pe_doing(pe_doing[13][5]),
        .c1_vld(c1_vld[13][5]),
        .c1_data(c1_data[13][47:40])
    );
    
    pe u_pe_row13_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[6]),
        .in0_data(sys_arr_row13_data[55:48]),
        .in1_vld(sys_arr_col6_vld[13]),
        .in1_data(sys_arr_col6_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[6]),
        .out0_data(sys_arr_row14_data[55:48]),
        .out1_vld(sys_arr_col7_vld[13]),
        .out1_data(sys_arr_col7_data[111:104]),
        .pe_doing(pe_doing[13][6]),
        .c1_vld(c1_vld[13][6]),
        .c1_data(c1_data[13][55:48])
    );
    
    pe u_pe_row13_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[7]),
        .in0_data(sys_arr_row13_data[63:56]),
        .in1_vld(sys_arr_col7_vld[13]),
        .in1_data(sys_arr_col7_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[7]),
        .out0_data(sys_arr_row14_data[63:56]),
        .out1_vld(sys_arr_col8_vld[13]),
        .out1_data(sys_arr_col8_data[111:104]),
        .pe_doing(pe_doing[13][7]),
        .c1_vld(c1_vld[13][7]),
        .c1_data(c1_data[13][63:56])
    );
    
    pe u_pe_row13_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[8]),
        .in0_data(sys_arr_row13_data[71:64]),
        .in1_vld(sys_arr_col8_vld[13]),
        .in1_data(sys_arr_col8_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[8]),
        .out0_data(sys_arr_row14_data[71:64]),
        .out1_vld(sys_arr_col9_vld[13]),
        .out1_data(sys_arr_col9_data[111:104]),
        .pe_doing(pe_doing[13][8]),
        .c1_vld(c1_vld[13][8]),
        .c1_data(c1_data[13][71:64])
    );
    
    pe u_pe_row13_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[9]),
        .in0_data(sys_arr_row13_data[79:72]),
        .in1_vld(sys_arr_col9_vld[13]),
        .in1_data(sys_arr_col9_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[9]),
        .out0_data(sys_arr_row14_data[79:72]),
        .out1_vld(sys_arr_col10_vld[13]),
        .out1_data(sys_arr_col10_data[111:104]),
        .pe_doing(pe_doing[13][9]),
        .c1_vld(c1_vld[13][9]),
        .c1_data(c1_data[13][79:72])
    );
    
    pe u_pe_row13_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[10]),
        .in0_data(sys_arr_row13_data[87:80]),
        .in1_vld(sys_arr_col10_vld[13]),
        .in1_data(sys_arr_col10_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[10]),
        .out0_data(sys_arr_row14_data[87:80]),
        .out1_vld(sys_arr_col11_vld[13]),
        .out1_data(sys_arr_col11_data[111:104]),
        .pe_doing(pe_doing[13][10]),
        .c1_vld(c1_vld[13][10]),
        .c1_data(c1_data[13][87:80])
    );
    
    pe u_pe_row13_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[11]),
        .in0_data(sys_arr_row13_data[95:88]),
        .in1_vld(sys_arr_col11_vld[13]),
        .in1_data(sys_arr_col11_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[11]),
        .out0_data(sys_arr_row14_data[95:88]),
        .out1_vld(sys_arr_col12_vld[13]),
        .out1_data(sys_arr_col12_data[111:104]),
        .pe_doing(pe_doing[13][11]),
        .c1_vld(c1_vld[13][11]),
        .c1_data(c1_data[13][95:88])
    );
    
    pe u_pe_row13_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[12]),
        .in0_data(sys_arr_row13_data[103:96]),
        .in1_vld(sys_arr_col12_vld[13]),
        .in1_data(sys_arr_col12_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[12]),
        .out0_data(sys_arr_row14_data[103:96]),
        .out1_vld(sys_arr_col13_vld[13]),
        .out1_data(sys_arr_col13_data[111:104]),
        .pe_doing(pe_doing[13][12]),
        .c1_vld(c1_vld[13][12]),
        .c1_data(c1_data[13][103:96])
    );
    
    pe u_pe_row13_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[13]),
        .in0_data(sys_arr_row13_data[111:104]),
        .in1_vld(sys_arr_col13_vld[13]),
        .in1_data(sys_arr_col13_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[13]),
        .out0_data(sys_arr_row14_data[111:104]),
        .out1_vld(sys_arr_col14_vld[13]),
        .out1_data(sys_arr_col14_data[111:104]),
        .pe_doing(pe_doing[13][13]),
        .c1_vld(c1_vld[13][13]),
        .c1_data(c1_data[13][111:104])
    );
    
    pe u_pe_row13_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[14]),
        .in0_data(sys_arr_row13_data[119:112]),
        .in1_vld(sys_arr_col14_vld[13]),
        .in1_data(sys_arr_col14_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[14]),
        .out0_data(sys_arr_row14_data[119:112]),
        .out1_vld(sys_arr_col15_vld[13]),
        .out1_data(sys_arr_col15_data[111:104]),
        .pe_doing(pe_doing[13][14]),
        .c1_vld(c1_vld[13][14]),
        .c1_data(c1_data[13][119:112])
    );
    
    pe u_pe_row13_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row13_vld[15]),
        .in0_data(sys_arr_row13_data[127:120]),
        .in1_vld(sys_arr_col15_vld[13]),
        .in1_data(sys_arr_col15_data[111:104]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row14_vld[15]),
        .out0_data(sys_arr_row14_data[127:120]),
        .out1_vld(sys_arr_col16_vld[13]),
        .out1_data(sys_arr_col16_data[111:104]),
        .pe_doing(pe_doing[13][15]),
        .c1_vld(c1_vld[13][15]),
        .c1_data(c1_data[13][127:120])
    );
    
    pe u_pe_row14_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[0]),
        .in0_data(sys_arr_row14_data[7:0]),
        .in1_vld(sys_arr_col0_vld[14]),
        .in1_data(sys_arr_col0_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[0]),
        .out0_data(sys_arr_row15_data[7:0]),
        .out1_vld(sys_arr_col1_vld[14]),
        .out1_data(sys_arr_col1_data[119:112]),
        .pe_doing(pe_doing[14][0]),
        .c1_vld(c1_vld[14][0]),
        .c1_data(c1_data[14][7:0])
    );
    
    pe u_pe_row14_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[1]),
        .in0_data(sys_arr_row14_data[15:8]),
        .in1_vld(sys_arr_col1_vld[14]),
        .in1_data(sys_arr_col1_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[1]),
        .out0_data(sys_arr_row15_data[15:8]),
        .out1_vld(sys_arr_col2_vld[14]),
        .out1_data(sys_arr_col2_data[119:112]),
        .pe_doing(pe_doing[14][1]),
        .c1_vld(c1_vld[14][1]),
        .c1_data(c1_data[14][15:8])
    );
    
    pe u_pe_row14_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[2]),
        .in0_data(sys_arr_row14_data[23:16]),
        .in1_vld(sys_arr_col2_vld[14]),
        .in1_data(sys_arr_col2_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[2]),
        .out0_data(sys_arr_row15_data[23:16]),
        .out1_vld(sys_arr_col3_vld[14]),
        .out1_data(sys_arr_col3_data[119:112]),
        .pe_doing(pe_doing[14][2]),
        .c1_vld(c1_vld[14][2]),
        .c1_data(c1_data[14][23:16])
    );
    
    pe u_pe_row14_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[3]),
        .in0_data(sys_arr_row14_data[31:24]),
        .in1_vld(sys_arr_col3_vld[14]),
        .in1_data(sys_arr_col3_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[3]),
        .out0_data(sys_arr_row15_data[31:24]),
        .out1_vld(sys_arr_col4_vld[14]),
        .out1_data(sys_arr_col4_data[119:112]),
        .pe_doing(pe_doing[14][3]),
        .c1_vld(c1_vld[14][3]),
        .c1_data(c1_data[14][31:24])
    );
    
    pe u_pe_row14_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[4]),
        .in0_data(sys_arr_row14_data[39:32]),
        .in1_vld(sys_arr_col4_vld[14]),
        .in1_data(sys_arr_col4_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[4]),
        .out0_data(sys_arr_row15_data[39:32]),
        .out1_vld(sys_arr_col5_vld[14]),
        .out1_data(sys_arr_col5_data[119:112]),
        .pe_doing(pe_doing[14][4]),
        .c1_vld(c1_vld[14][4]),
        .c1_data(c1_data[14][39:32])
    );
    
    pe u_pe_row14_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[5]),
        .in0_data(sys_arr_row14_data[47:40]),
        .in1_vld(sys_arr_col5_vld[14]),
        .in1_data(sys_arr_col5_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[5]),
        .out0_data(sys_arr_row15_data[47:40]),
        .out1_vld(sys_arr_col6_vld[14]),
        .out1_data(sys_arr_col6_data[119:112]),
        .pe_doing(pe_doing[14][5]),
        .c1_vld(c1_vld[14][5]),
        .c1_data(c1_data[14][47:40])
    );
    
    pe u_pe_row14_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[6]),
        .in0_data(sys_arr_row14_data[55:48]),
        .in1_vld(sys_arr_col6_vld[14]),
        .in1_data(sys_arr_col6_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[6]),
        .out0_data(sys_arr_row15_data[55:48]),
        .out1_vld(sys_arr_col7_vld[14]),
        .out1_data(sys_arr_col7_data[119:112]),
        .pe_doing(pe_doing[14][6]),
        .c1_vld(c1_vld[14][6]),
        .c1_data(c1_data[14][55:48])
    );
    
    pe u_pe_row14_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[7]),
        .in0_data(sys_arr_row14_data[63:56]),
        .in1_vld(sys_arr_col7_vld[14]),
        .in1_data(sys_arr_col7_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[7]),
        .out0_data(sys_arr_row15_data[63:56]),
        .out1_vld(sys_arr_col8_vld[14]),
        .out1_data(sys_arr_col8_data[119:112]),
        .pe_doing(pe_doing[14][7]),
        .c1_vld(c1_vld[14][7]),
        .c1_data(c1_data[14][63:56])
    );
    
    pe u_pe_row14_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[8]),
        .in0_data(sys_arr_row14_data[71:64]),
        .in1_vld(sys_arr_col8_vld[14]),
        .in1_data(sys_arr_col8_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[8]),
        .out0_data(sys_arr_row15_data[71:64]),
        .out1_vld(sys_arr_col9_vld[14]),
        .out1_data(sys_arr_col9_data[119:112]),
        .pe_doing(pe_doing[14][8]),
        .c1_vld(c1_vld[14][8]),
        .c1_data(c1_data[14][71:64])
    );
    
    pe u_pe_row14_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[9]),
        .in0_data(sys_arr_row14_data[79:72]),
        .in1_vld(sys_arr_col9_vld[14]),
        .in1_data(sys_arr_col9_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[9]),
        .out0_data(sys_arr_row15_data[79:72]),
        .out1_vld(sys_arr_col10_vld[14]),
        .out1_data(sys_arr_col10_data[119:112]),
        .pe_doing(pe_doing[14][9]),
        .c1_vld(c1_vld[14][9]),
        .c1_data(c1_data[14][79:72])
    );
    
    pe u_pe_row14_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[10]),
        .in0_data(sys_arr_row14_data[87:80]),
        .in1_vld(sys_arr_col10_vld[14]),
        .in1_data(sys_arr_col10_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[10]),
        .out0_data(sys_arr_row15_data[87:80]),
        .out1_vld(sys_arr_col11_vld[14]),
        .out1_data(sys_arr_col11_data[119:112]),
        .pe_doing(pe_doing[14][10]),
        .c1_vld(c1_vld[14][10]),
        .c1_data(c1_data[14][87:80])
    );
    
    pe u_pe_row14_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[11]),
        .in0_data(sys_arr_row14_data[95:88]),
        .in1_vld(sys_arr_col11_vld[14]),
        .in1_data(sys_arr_col11_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[11]),
        .out0_data(sys_arr_row15_data[95:88]),
        .out1_vld(sys_arr_col12_vld[14]),
        .out1_data(sys_arr_col12_data[119:112]),
        .pe_doing(pe_doing[14][11]),
        .c1_vld(c1_vld[14][11]),
        .c1_data(c1_data[14][95:88])
    );
    
    pe u_pe_row14_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[12]),
        .in0_data(sys_arr_row14_data[103:96]),
        .in1_vld(sys_arr_col12_vld[14]),
        .in1_data(sys_arr_col12_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[12]),
        .out0_data(sys_arr_row15_data[103:96]),
        .out1_vld(sys_arr_col13_vld[14]),
        .out1_data(sys_arr_col13_data[119:112]),
        .pe_doing(pe_doing[14][12]),
        .c1_vld(c1_vld[14][12]),
        .c1_data(c1_data[14][103:96])
    );
    
    pe u_pe_row14_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[13]),
        .in0_data(sys_arr_row14_data[111:104]),
        .in1_vld(sys_arr_col13_vld[14]),
        .in1_data(sys_arr_col13_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[13]),
        .out0_data(sys_arr_row15_data[111:104]),
        .out1_vld(sys_arr_col14_vld[14]),
        .out1_data(sys_arr_col14_data[119:112]),
        .pe_doing(pe_doing[14][13]),
        .c1_vld(c1_vld[14][13]),
        .c1_data(c1_data[14][111:104])
    );
    
    pe u_pe_row14_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[14]),
        .in0_data(sys_arr_row14_data[119:112]),
        .in1_vld(sys_arr_col14_vld[14]),
        .in1_data(sys_arr_col14_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[14]),
        .out0_data(sys_arr_row15_data[119:112]),
        .out1_vld(sys_arr_col15_vld[14]),
        .out1_data(sys_arr_col15_data[119:112]),
        .pe_doing(pe_doing[14][14]),
        .c1_vld(c1_vld[14][14]),
        .c1_data(c1_data[14][119:112])
    );
    
    pe u_pe_row14_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row14_vld[15]),
        .in0_data(sys_arr_row14_data[127:120]),
        .in1_vld(sys_arr_col15_vld[14]),
        .in1_data(sys_arr_col15_data[119:112]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row15_vld[15]),
        .out0_data(sys_arr_row15_data[127:120]),
        .out1_vld(sys_arr_col16_vld[14]),
        .out1_data(sys_arr_col16_data[119:112]),
        .pe_doing(pe_doing[14][15]),
        .c1_vld(c1_vld[14][15]),
        .c1_data(c1_data[14][127:120])
    );
    
    pe u_pe_row15_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[0]),
        .in0_data(sys_arr_row15_data[7:0]),
        .in1_vld(sys_arr_col0_vld[15]),
        .in1_data(sys_arr_col0_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[0]),
        .out0_data(sys_arr_row16_data[7:0]),
        .out1_vld(sys_arr_col1_vld[15]),
        .out1_data(sys_arr_col1_data[127:120]),
        .pe_doing(pe_doing[15][0]),
        .c1_vld(c1_vld[15][0]),
        .c1_data(c1_data[15][7:0])
    );
    
    pe u_pe_row15_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[1]),
        .in0_data(sys_arr_row15_data[15:8]),
        .in1_vld(sys_arr_col1_vld[15]),
        .in1_data(sys_arr_col1_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[1]),
        .out0_data(sys_arr_row16_data[15:8]),
        .out1_vld(sys_arr_col2_vld[15]),
        .out1_data(sys_arr_col2_data[127:120]),
        .pe_doing(pe_doing[15][1]),
        .c1_vld(c1_vld[15][1]),
        .c1_data(c1_data[15][15:8])
    );
    
    pe u_pe_row15_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[2]),
        .in0_data(sys_arr_row15_data[23:16]),
        .in1_vld(sys_arr_col2_vld[15]),
        .in1_data(sys_arr_col2_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[2]),
        .out0_data(sys_arr_row16_data[23:16]),
        .out1_vld(sys_arr_col3_vld[15]),
        .out1_data(sys_arr_col3_data[127:120]),
        .pe_doing(pe_doing[15][2]),
        .c1_vld(c1_vld[15][2]),
        .c1_data(c1_data[15][23:16])
    );
    
    pe u_pe_row15_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[3]),
        .in0_data(sys_arr_row15_data[31:24]),
        .in1_vld(sys_arr_col3_vld[15]),
        .in1_data(sys_arr_col3_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[3]),
        .out0_data(sys_arr_row16_data[31:24]),
        .out1_vld(sys_arr_col4_vld[15]),
        .out1_data(sys_arr_col4_data[127:120]),
        .pe_doing(pe_doing[15][3]),
        .c1_vld(c1_vld[15][3]),
        .c1_data(c1_data[15][31:24])
    );
    
    pe u_pe_row15_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[4]),
        .in0_data(sys_arr_row15_data[39:32]),
        .in1_vld(sys_arr_col4_vld[15]),
        .in1_data(sys_arr_col4_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[4]),
        .out0_data(sys_arr_row16_data[39:32]),
        .out1_vld(sys_arr_col5_vld[15]),
        .out1_data(sys_arr_col5_data[127:120]),
        .pe_doing(pe_doing[15][4]),
        .c1_vld(c1_vld[15][4]),
        .c1_data(c1_data[15][39:32])
    );
    
    pe u_pe_row15_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[5]),
        .in0_data(sys_arr_row15_data[47:40]),
        .in1_vld(sys_arr_col5_vld[15]),
        .in1_data(sys_arr_col5_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[5]),
        .out0_data(sys_arr_row16_data[47:40]),
        .out1_vld(sys_arr_col6_vld[15]),
        .out1_data(sys_arr_col6_data[127:120]),
        .pe_doing(pe_doing[15][5]),
        .c1_vld(c1_vld[15][5]),
        .c1_data(c1_data[15][47:40])
    );
    
    pe u_pe_row15_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[6]),
        .in0_data(sys_arr_row15_data[55:48]),
        .in1_vld(sys_arr_col6_vld[15]),
        .in1_data(sys_arr_col6_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[6]),
        .out0_data(sys_arr_row16_data[55:48]),
        .out1_vld(sys_arr_col7_vld[15]),
        .out1_data(sys_arr_col7_data[127:120]),
        .pe_doing(pe_doing[15][6]),
        .c1_vld(c1_vld[15][6]),
        .c1_data(c1_data[15][55:48])
    );
    
    pe u_pe_row15_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[7]),
        .in0_data(sys_arr_row15_data[63:56]),
        .in1_vld(sys_arr_col7_vld[15]),
        .in1_data(sys_arr_col7_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[7]),
        .out0_data(sys_arr_row16_data[63:56]),
        .out1_vld(sys_arr_col8_vld[15]),
        .out1_data(sys_arr_col8_data[127:120]),
        .pe_doing(pe_doing[15][7]),
        .c1_vld(c1_vld[15][7]),
        .c1_data(c1_data[15][63:56])
    );
    
    pe u_pe_row15_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[8]),
        .in0_data(sys_arr_row15_data[71:64]),
        .in1_vld(sys_arr_col8_vld[15]),
        .in1_data(sys_arr_col8_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[8]),
        .out0_data(sys_arr_row16_data[71:64]),
        .out1_vld(sys_arr_col9_vld[15]),
        .out1_data(sys_arr_col9_data[127:120]),
        .pe_doing(pe_doing[15][8]),
        .c1_vld(c1_vld[15][8]),
        .c1_data(c1_data[15][71:64])
    );
    
    pe u_pe_row15_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[9]),
        .in0_data(sys_arr_row15_data[79:72]),
        .in1_vld(sys_arr_col9_vld[15]),
        .in1_data(sys_arr_col9_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[9]),
        .out0_data(sys_arr_row16_data[79:72]),
        .out1_vld(sys_arr_col10_vld[15]),
        .out1_data(sys_arr_col10_data[127:120]),
        .pe_doing(pe_doing[15][9]),
        .c1_vld(c1_vld[15][9]),
        .c1_data(c1_data[15][79:72])
    );
    
    pe u_pe_row15_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[10]),
        .in0_data(sys_arr_row15_data[87:80]),
        .in1_vld(sys_arr_col10_vld[15]),
        .in1_data(sys_arr_col10_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[10]),
        .out0_data(sys_arr_row16_data[87:80]),
        .out1_vld(sys_arr_col11_vld[15]),
        .out1_data(sys_arr_col11_data[127:120]),
        .pe_doing(pe_doing[15][10]),
        .c1_vld(c1_vld[15][10]),
        .c1_data(c1_data[15][87:80])
    );
    
    pe u_pe_row15_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[11]),
        .in0_data(sys_arr_row15_data[95:88]),
        .in1_vld(sys_arr_col11_vld[15]),
        .in1_data(sys_arr_col11_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[11]),
        .out0_data(sys_arr_row16_data[95:88]),
        .out1_vld(sys_arr_col12_vld[15]),
        .out1_data(sys_arr_col12_data[127:120]),
        .pe_doing(pe_doing[15][11]),
        .c1_vld(c1_vld[15][11]),
        .c1_data(c1_data[15][95:88])
    );
    
    pe u_pe_row15_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[12]),
        .in0_data(sys_arr_row15_data[103:96]),
        .in1_vld(sys_arr_col12_vld[15]),
        .in1_data(sys_arr_col12_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[12]),
        .out0_data(sys_arr_row16_data[103:96]),
        .out1_vld(sys_arr_col13_vld[15]),
        .out1_data(sys_arr_col13_data[127:120]),
        .pe_doing(pe_doing[15][12]),
        .c1_vld(c1_vld[15][12]),
        .c1_data(c1_data[15][103:96])
    );
    
    pe u_pe_row15_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[13]),
        .in0_data(sys_arr_row15_data[111:104]),
        .in1_vld(sys_arr_col13_vld[15]),
        .in1_data(sys_arr_col13_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[13]),
        .out0_data(sys_arr_row16_data[111:104]),
        .out1_vld(sys_arr_col14_vld[15]),
        .out1_data(sys_arr_col14_data[127:120]),
        .pe_doing(pe_doing[15][13]),
        .c1_vld(c1_vld[15][13]),
        .c1_data(c1_data[15][111:104])
    );
    
    pe u_pe_row15_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[14]),
        .in0_data(sys_arr_row15_data[119:112]),
        .in1_vld(sys_arr_col14_vld[15]),
        .in1_data(sys_arr_col14_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[14]),
        .out0_data(sys_arr_row16_data[119:112]),
        .out1_vld(sys_arr_col15_vld[15]),
        .out1_data(sys_arr_col15_data[127:120]),
        .pe_doing(pe_doing[15][14]),
        .c1_vld(c1_vld[15][14]),
        .c1_data(c1_data[15][119:112])
    );
    
    pe u_pe_row15_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .in0_vld(sys_arr_row15_vld[15]),
        .in0_data(sys_arr_row15_data[127:120]),
        .in1_vld(sys_arr_col15_vld[15]),
        .in1_data(sys_arr_col15_data[127:120]),
        .pe_en(mxu_vld),
        .out0_vld(sys_arr_row16_vld[15]),
        .out0_data(sys_arr_row16_data[127:120]),
        .out1_vld(sys_arr_col16_vld[15]),
        .out1_data(sys_arr_col16_data[127:120]),
        .pe_doing(pe_doing[15][15]),
        .c1_vld(c1_vld[15][15]),
        .c1_data(c1_data[15][127:120])
    );
    

    acc u_acc_row0_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][0]),
        .acc_data(c1_data[0][7:0]),
        .load_vld(sys_arr_row0_load_vld[0]),
        .load_data(sys_arr_row0_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row0_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row0_data[7:0])
    );
    
    acc u_acc_row0_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][1]),
        .acc_data(c1_data[0][15:8]),
        .load_vld(sys_arr_row0_load_vld[1]),
        .load_data(sys_arr_row0_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row0_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row0_data[15:8])
    );
    
    acc u_acc_row0_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][2]),
        .acc_data(c1_data[0][23:16]),
        .load_vld(sys_arr_row0_load_vld[2]),
        .load_data(sys_arr_row0_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row0_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row0_data[23:16])
    );
    
    acc u_acc_row0_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][3]),
        .acc_data(c1_data[0][31:24]),
        .load_vld(sys_arr_row0_load_vld[3]),
        .load_data(sys_arr_row0_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row0_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row0_data[31:24])
    );
    
    acc u_acc_row0_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][4]),
        .acc_data(c1_data[0][39:32]),
        .load_vld(sys_arr_row0_load_vld[4]),
        .load_data(sys_arr_row0_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row0_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row0_data[39:32])
    );
    
    acc u_acc_row0_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][5]),
        .acc_data(c1_data[0][47:40]),
        .load_vld(sys_arr_row0_load_vld[5]),
        .load_data(sys_arr_row0_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row0_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row0_data[47:40])
    );
    
    acc u_acc_row0_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][6]),
        .acc_data(c1_data[0][55:48]),
        .load_vld(sys_arr_row0_load_vld[6]),
        .load_data(sys_arr_row0_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row0_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row0_data[55:48])
    );
    
    acc u_acc_row0_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][7]),
        .acc_data(c1_data[0][63:56]),
        .load_vld(sys_arr_row0_load_vld[7]),
        .load_data(sys_arr_row0_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row0_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row0_data[63:56])
    );
    
    acc u_acc_row0_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][8]),
        .acc_data(c1_data[0][71:64]),
        .load_vld(sys_arr_row0_load_vld[8]),
        .load_data(sys_arr_row0_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row0_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row0_data[71:64])
    );
    
    acc u_acc_row0_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][9]),
        .acc_data(c1_data[0][79:72]),
        .load_vld(sys_arr_row0_load_vld[9]),
        .load_data(sys_arr_row0_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row0_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row0_data[79:72])
    );
    
    acc u_acc_row0_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][10]),
        .acc_data(c1_data[0][87:80]),
        .load_vld(sys_arr_row0_load_vld[10]),
        .load_data(sys_arr_row0_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row0_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row0_data[87:80])
    );
    
    acc u_acc_row0_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][11]),
        .acc_data(c1_data[0][95:88]),
        .load_vld(sys_arr_row0_load_vld[11]),
        .load_data(sys_arr_row0_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row0_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row0_data[95:88])
    );
    
    acc u_acc_row0_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][12]),
        .acc_data(c1_data[0][103:96]),
        .load_vld(sys_arr_row0_load_vld[12]),
        .load_data(sys_arr_row0_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row0_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row0_data[103:96])
    );
    
    acc u_acc_row0_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][13]),
        .acc_data(c1_data[0][111:104]),
        .load_vld(sys_arr_row0_load_vld[13]),
        .load_data(sys_arr_row0_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row0_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row0_data[111:104])
    );
    
    acc u_acc_row0_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][14]),
        .acc_data(c1_data[0][119:112]),
        .load_vld(sys_arr_row0_load_vld[14]),
        .load_data(sys_arr_row0_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row0_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row0_data[119:112])
    );
    
    acc u_acc_row0_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[0][15]),
        .acc_data(c1_data[0][127:120]),
        .load_vld(sys_arr_row0_load_vld[15]),
        .load_data(sys_arr_row0_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row0_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row0_data[127:120])
    );
    
    acc u_acc_row1_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][0]),
        .acc_data(c1_data[1][7:0]),
        .load_vld(sys_arr_row1_load_vld[0]),
        .load_data(sys_arr_row1_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row1_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row1_data[7:0])
    );
    
    acc u_acc_row1_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][1]),
        .acc_data(c1_data[1][15:8]),
        .load_vld(sys_arr_row1_load_vld[1]),
        .load_data(sys_arr_row1_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row1_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row1_data[15:8])
    );
    
    acc u_acc_row1_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][2]),
        .acc_data(c1_data[1][23:16]),
        .load_vld(sys_arr_row1_load_vld[2]),
        .load_data(sys_arr_row1_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row1_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row1_data[23:16])
    );
    
    acc u_acc_row1_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][3]),
        .acc_data(c1_data[1][31:24]),
        .load_vld(sys_arr_row1_load_vld[3]),
        .load_data(sys_arr_row1_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row1_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row1_data[31:24])
    );
    
    acc u_acc_row1_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][4]),
        .acc_data(c1_data[1][39:32]),
        .load_vld(sys_arr_row1_load_vld[4]),
        .load_data(sys_arr_row1_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row1_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row1_data[39:32])
    );
    
    acc u_acc_row1_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][5]),
        .acc_data(c1_data[1][47:40]),
        .load_vld(sys_arr_row1_load_vld[5]),
        .load_data(sys_arr_row1_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row1_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row1_data[47:40])
    );
    
    acc u_acc_row1_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][6]),
        .acc_data(c1_data[1][55:48]),
        .load_vld(sys_arr_row1_load_vld[6]),
        .load_data(sys_arr_row1_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row1_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row1_data[55:48])
    );
    
    acc u_acc_row1_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][7]),
        .acc_data(c1_data[1][63:56]),
        .load_vld(sys_arr_row1_load_vld[7]),
        .load_data(sys_arr_row1_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row1_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row1_data[63:56])
    );
    
    acc u_acc_row1_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][8]),
        .acc_data(c1_data[1][71:64]),
        .load_vld(sys_arr_row1_load_vld[8]),
        .load_data(sys_arr_row1_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row1_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row1_data[71:64])
    );
    
    acc u_acc_row1_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][9]),
        .acc_data(c1_data[1][79:72]),
        .load_vld(sys_arr_row1_load_vld[9]),
        .load_data(sys_arr_row1_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row1_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row1_data[79:72])
    );
    
    acc u_acc_row1_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][10]),
        .acc_data(c1_data[1][87:80]),
        .load_vld(sys_arr_row1_load_vld[10]),
        .load_data(sys_arr_row1_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row1_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row1_data[87:80])
    );
    
    acc u_acc_row1_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][11]),
        .acc_data(c1_data[1][95:88]),
        .load_vld(sys_arr_row1_load_vld[11]),
        .load_data(sys_arr_row1_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row1_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row1_data[95:88])
    );
    
    acc u_acc_row1_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][12]),
        .acc_data(c1_data[1][103:96]),
        .load_vld(sys_arr_row1_load_vld[12]),
        .load_data(sys_arr_row1_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row1_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row1_data[103:96])
    );
    
    acc u_acc_row1_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][13]),
        .acc_data(c1_data[1][111:104]),
        .load_vld(sys_arr_row1_load_vld[13]),
        .load_data(sys_arr_row1_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row1_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row1_data[111:104])
    );
    
    acc u_acc_row1_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][14]),
        .acc_data(c1_data[1][119:112]),
        .load_vld(sys_arr_row1_load_vld[14]),
        .load_data(sys_arr_row1_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row1_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row1_data[119:112])
    );
    
    acc u_acc_row1_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[1][15]),
        .acc_data(c1_data[1][127:120]),
        .load_vld(sys_arr_row1_load_vld[15]),
        .load_data(sys_arr_row1_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row1_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row1_data[127:120])
    );
    
    acc u_acc_row2_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][0]),
        .acc_data(c1_data[2][7:0]),
        .load_vld(sys_arr_row2_load_vld[0]),
        .load_data(sys_arr_row2_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row2_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row2_data[7:0])
    );
    
    acc u_acc_row2_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][1]),
        .acc_data(c1_data[2][15:8]),
        .load_vld(sys_arr_row2_load_vld[1]),
        .load_data(sys_arr_row2_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row2_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row2_data[15:8])
    );
    
    acc u_acc_row2_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][2]),
        .acc_data(c1_data[2][23:16]),
        .load_vld(sys_arr_row2_load_vld[2]),
        .load_data(sys_arr_row2_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row2_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row2_data[23:16])
    );
    
    acc u_acc_row2_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][3]),
        .acc_data(c1_data[2][31:24]),
        .load_vld(sys_arr_row2_load_vld[3]),
        .load_data(sys_arr_row2_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row2_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row2_data[31:24])
    );
    
    acc u_acc_row2_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][4]),
        .acc_data(c1_data[2][39:32]),
        .load_vld(sys_arr_row2_load_vld[4]),
        .load_data(sys_arr_row2_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row2_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row2_data[39:32])
    );
    
    acc u_acc_row2_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][5]),
        .acc_data(c1_data[2][47:40]),
        .load_vld(sys_arr_row2_load_vld[5]),
        .load_data(sys_arr_row2_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row2_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row2_data[47:40])
    );
    
    acc u_acc_row2_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][6]),
        .acc_data(c1_data[2][55:48]),
        .load_vld(sys_arr_row2_load_vld[6]),
        .load_data(sys_arr_row2_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row2_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row2_data[55:48])
    );
    
    acc u_acc_row2_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][7]),
        .acc_data(c1_data[2][63:56]),
        .load_vld(sys_arr_row2_load_vld[7]),
        .load_data(sys_arr_row2_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row2_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row2_data[63:56])
    );
    
    acc u_acc_row2_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][8]),
        .acc_data(c1_data[2][71:64]),
        .load_vld(sys_arr_row2_load_vld[8]),
        .load_data(sys_arr_row2_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row2_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row2_data[71:64])
    );
    
    acc u_acc_row2_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][9]),
        .acc_data(c1_data[2][79:72]),
        .load_vld(sys_arr_row2_load_vld[9]),
        .load_data(sys_arr_row2_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row2_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row2_data[79:72])
    );
    
    acc u_acc_row2_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][10]),
        .acc_data(c1_data[2][87:80]),
        .load_vld(sys_arr_row2_load_vld[10]),
        .load_data(sys_arr_row2_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row2_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row2_data[87:80])
    );
    
    acc u_acc_row2_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][11]),
        .acc_data(c1_data[2][95:88]),
        .load_vld(sys_arr_row2_load_vld[11]),
        .load_data(sys_arr_row2_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row2_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row2_data[95:88])
    );
    
    acc u_acc_row2_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][12]),
        .acc_data(c1_data[2][103:96]),
        .load_vld(sys_arr_row2_load_vld[12]),
        .load_data(sys_arr_row2_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row2_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row2_data[103:96])
    );
    
    acc u_acc_row2_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][13]),
        .acc_data(c1_data[2][111:104]),
        .load_vld(sys_arr_row2_load_vld[13]),
        .load_data(sys_arr_row2_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row2_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row2_data[111:104])
    );
    
    acc u_acc_row2_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][14]),
        .acc_data(c1_data[2][119:112]),
        .load_vld(sys_arr_row2_load_vld[14]),
        .load_data(sys_arr_row2_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row2_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row2_data[119:112])
    );
    
    acc u_acc_row2_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[2][15]),
        .acc_data(c1_data[2][127:120]),
        .load_vld(sys_arr_row2_load_vld[15]),
        .load_data(sys_arr_row2_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row2_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row2_data[127:120])
    );
    
    acc u_acc_row3_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][0]),
        .acc_data(c1_data[3][7:0]),
        .load_vld(sys_arr_row3_load_vld[0]),
        .load_data(sys_arr_row3_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row3_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row3_data[7:0])
    );
    
    acc u_acc_row3_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][1]),
        .acc_data(c1_data[3][15:8]),
        .load_vld(sys_arr_row3_load_vld[1]),
        .load_data(sys_arr_row3_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row3_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row3_data[15:8])
    );
    
    acc u_acc_row3_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][2]),
        .acc_data(c1_data[3][23:16]),
        .load_vld(sys_arr_row3_load_vld[2]),
        .load_data(sys_arr_row3_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row3_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row3_data[23:16])
    );
    
    acc u_acc_row3_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][3]),
        .acc_data(c1_data[3][31:24]),
        .load_vld(sys_arr_row3_load_vld[3]),
        .load_data(sys_arr_row3_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row3_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row3_data[31:24])
    );
    
    acc u_acc_row3_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][4]),
        .acc_data(c1_data[3][39:32]),
        .load_vld(sys_arr_row3_load_vld[4]),
        .load_data(sys_arr_row3_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row3_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row3_data[39:32])
    );
    
    acc u_acc_row3_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][5]),
        .acc_data(c1_data[3][47:40]),
        .load_vld(sys_arr_row3_load_vld[5]),
        .load_data(sys_arr_row3_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row3_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row3_data[47:40])
    );
    
    acc u_acc_row3_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][6]),
        .acc_data(c1_data[3][55:48]),
        .load_vld(sys_arr_row3_load_vld[6]),
        .load_data(sys_arr_row3_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row3_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row3_data[55:48])
    );
    
    acc u_acc_row3_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][7]),
        .acc_data(c1_data[3][63:56]),
        .load_vld(sys_arr_row3_load_vld[7]),
        .load_data(sys_arr_row3_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row3_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row3_data[63:56])
    );
    
    acc u_acc_row3_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][8]),
        .acc_data(c1_data[3][71:64]),
        .load_vld(sys_arr_row3_load_vld[8]),
        .load_data(sys_arr_row3_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row3_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row3_data[71:64])
    );
    
    acc u_acc_row3_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][9]),
        .acc_data(c1_data[3][79:72]),
        .load_vld(sys_arr_row3_load_vld[9]),
        .load_data(sys_arr_row3_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row3_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row3_data[79:72])
    );
    
    acc u_acc_row3_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][10]),
        .acc_data(c1_data[3][87:80]),
        .load_vld(sys_arr_row3_load_vld[10]),
        .load_data(sys_arr_row3_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row3_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row3_data[87:80])
    );
    
    acc u_acc_row3_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][11]),
        .acc_data(c1_data[3][95:88]),
        .load_vld(sys_arr_row3_load_vld[11]),
        .load_data(sys_arr_row3_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row3_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row3_data[95:88])
    );
    
    acc u_acc_row3_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][12]),
        .acc_data(c1_data[3][103:96]),
        .load_vld(sys_arr_row3_load_vld[12]),
        .load_data(sys_arr_row3_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row3_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row3_data[103:96])
    );
    
    acc u_acc_row3_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][13]),
        .acc_data(c1_data[3][111:104]),
        .load_vld(sys_arr_row3_load_vld[13]),
        .load_data(sys_arr_row3_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row3_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row3_data[111:104])
    );
    
    acc u_acc_row3_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][14]),
        .acc_data(c1_data[3][119:112]),
        .load_vld(sys_arr_row3_load_vld[14]),
        .load_data(sys_arr_row3_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row3_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row3_data[119:112])
    );
    
    acc u_acc_row3_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[3][15]),
        .acc_data(c1_data[3][127:120]),
        .load_vld(sys_arr_row3_load_vld[15]),
        .load_data(sys_arr_row3_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row3_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row3_data[127:120])
    );
    
    acc u_acc_row4_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][0]),
        .acc_data(c1_data[4][7:0]),
        .load_vld(sys_arr_row4_load_vld[0]),
        .load_data(sys_arr_row4_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row4_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row4_data[7:0])
    );
    
    acc u_acc_row4_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][1]),
        .acc_data(c1_data[4][15:8]),
        .load_vld(sys_arr_row4_load_vld[1]),
        .load_data(sys_arr_row4_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row4_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row4_data[15:8])
    );
    
    acc u_acc_row4_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][2]),
        .acc_data(c1_data[4][23:16]),
        .load_vld(sys_arr_row4_load_vld[2]),
        .load_data(sys_arr_row4_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row4_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row4_data[23:16])
    );
    
    acc u_acc_row4_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][3]),
        .acc_data(c1_data[4][31:24]),
        .load_vld(sys_arr_row4_load_vld[3]),
        .load_data(sys_arr_row4_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row4_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row4_data[31:24])
    );
    
    acc u_acc_row4_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][4]),
        .acc_data(c1_data[4][39:32]),
        .load_vld(sys_arr_row4_load_vld[4]),
        .load_data(sys_arr_row4_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row4_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row4_data[39:32])
    );
    
    acc u_acc_row4_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][5]),
        .acc_data(c1_data[4][47:40]),
        .load_vld(sys_arr_row4_load_vld[5]),
        .load_data(sys_arr_row4_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row4_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row4_data[47:40])
    );
    
    acc u_acc_row4_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][6]),
        .acc_data(c1_data[4][55:48]),
        .load_vld(sys_arr_row4_load_vld[6]),
        .load_data(sys_arr_row4_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row4_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row4_data[55:48])
    );
    
    acc u_acc_row4_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][7]),
        .acc_data(c1_data[4][63:56]),
        .load_vld(sys_arr_row4_load_vld[7]),
        .load_data(sys_arr_row4_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row4_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row4_data[63:56])
    );
    
    acc u_acc_row4_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][8]),
        .acc_data(c1_data[4][71:64]),
        .load_vld(sys_arr_row4_load_vld[8]),
        .load_data(sys_arr_row4_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row4_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row4_data[71:64])
    );
    
    acc u_acc_row4_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][9]),
        .acc_data(c1_data[4][79:72]),
        .load_vld(sys_arr_row4_load_vld[9]),
        .load_data(sys_arr_row4_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row4_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row4_data[79:72])
    );
    
    acc u_acc_row4_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][10]),
        .acc_data(c1_data[4][87:80]),
        .load_vld(sys_arr_row4_load_vld[10]),
        .load_data(sys_arr_row4_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row4_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row4_data[87:80])
    );
    
    acc u_acc_row4_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][11]),
        .acc_data(c1_data[4][95:88]),
        .load_vld(sys_arr_row4_load_vld[11]),
        .load_data(sys_arr_row4_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row4_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row4_data[95:88])
    );
    
    acc u_acc_row4_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][12]),
        .acc_data(c1_data[4][103:96]),
        .load_vld(sys_arr_row4_load_vld[12]),
        .load_data(sys_arr_row4_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row4_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row4_data[103:96])
    );
    
    acc u_acc_row4_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][13]),
        .acc_data(c1_data[4][111:104]),
        .load_vld(sys_arr_row4_load_vld[13]),
        .load_data(sys_arr_row4_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row4_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row4_data[111:104])
    );
    
    acc u_acc_row4_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][14]),
        .acc_data(c1_data[4][119:112]),
        .load_vld(sys_arr_row4_load_vld[14]),
        .load_data(sys_arr_row4_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row4_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row4_data[119:112])
    );
    
    acc u_acc_row4_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[4][15]),
        .acc_data(c1_data[4][127:120]),
        .load_vld(sys_arr_row4_load_vld[15]),
        .load_data(sys_arr_row4_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row4_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row4_data[127:120])
    );
    
    acc u_acc_row5_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][0]),
        .acc_data(c1_data[5][7:0]),
        .load_vld(sys_arr_row5_load_vld[0]),
        .load_data(sys_arr_row5_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row5_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row5_data[7:0])
    );
    
    acc u_acc_row5_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][1]),
        .acc_data(c1_data[5][15:8]),
        .load_vld(sys_arr_row5_load_vld[1]),
        .load_data(sys_arr_row5_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row5_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row5_data[15:8])
    );
    
    acc u_acc_row5_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][2]),
        .acc_data(c1_data[5][23:16]),
        .load_vld(sys_arr_row5_load_vld[2]),
        .load_data(sys_arr_row5_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row5_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row5_data[23:16])
    );
    
    acc u_acc_row5_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][3]),
        .acc_data(c1_data[5][31:24]),
        .load_vld(sys_arr_row5_load_vld[3]),
        .load_data(sys_arr_row5_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row5_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row5_data[31:24])
    );
    
    acc u_acc_row5_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][4]),
        .acc_data(c1_data[5][39:32]),
        .load_vld(sys_arr_row5_load_vld[4]),
        .load_data(sys_arr_row5_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row5_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row5_data[39:32])
    );
    
    acc u_acc_row5_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][5]),
        .acc_data(c1_data[5][47:40]),
        .load_vld(sys_arr_row5_load_vld[5]),
        .load_data(sys_arr_row5_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row5_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row5_data[47:40])
    );
    
    acc u_acc_row5_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][6]),
        .acc_data(c1_data[5][55:48]),
        .load_vld(sys_arr_row5_load_vld[6]),
        .load_data(sys_arr_row5_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row5_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row5_data[55:48])
    );
    
    acc u_acc_row5_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][7]),
        .acc_data(c1_data[5][63:56]),
        .load_vld(sys_arr_row5_load_vld[7]),
        .load_data(sys_arr_row5_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row5_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row5_data[63:56])
    );
    
    acc u_acc_row5_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][8]),
        .acc_data(c1_data[5][71:64]),
        .load_vld(sys_arr_row5_load_vld[8]),
        .load_data(sys_arr_row5_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row5_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row5_data[71:64])
    );
    
    acc u_acc_row5_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][9]),
        .acc_data(c1_data[5][79:72]),
        .load_vld(sys_arr_row5_load_vld[9]),
        .load_data(sys_arr_row5_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row5_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row5_data[79:72])
    );
    
    acc u_acc_row5_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][10]),
        .acc_data(c1_data[5][87:80]),
        .load_vld(sys_arr_row5_load_vld[10]),
        .load_data(sys_arr_row5_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row5_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row5_data[87:80])
    );
    
    acc u_acc_row5_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][11]),
        .acc_data(c1_data[5][95:88]),
        .load_vld(sys_arr_row5_load_vld[11]),
        .load_data(sys_arr_row5_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row5_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row5_data[95:88])
    );
    
    acc u_acc_row5_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][12]),
        .acc_data(c1_data[5][103:96]),
        .load_vld(sys_arr_row5_load_vld[12]),
        .load_data(sys_arr_row5_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row5_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row5_data[103:96])
    );
    
    acc u_acc_row5_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][13]),
        .acc_data(c1_data[5][111:104]),
        .load_vld(sys_arr_row5_load_vld[13]),
        .load_data(sys_arr_row5_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row5_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row5_data[111:104])
    );
    
    acc u_acc_row5_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][14]),
        .acc_data(c1_data[5][119:112]),
        .load_vld(sys_arr_row5_load_vld[14]),
        .load_data(sys_arr_row5_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row5_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row5_data[119:112])
    );
    
    acc u_acc_row5_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[5][15]),
        .acc_data(c1_data[5][127:120]),
        .load_vld(sys_arr_row5_load_vld[15]),
        .load_data(sys_arr_row5_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row5_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row5_data[127:120])
    );
    
    acc u_acc_row6_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][0]),
        .acc_data(c1_data[6][7:0]),
        .load_vld(sys_arr_row6_load_vld[0]),
        .load_data(sys_arr_row6_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row6_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row6_data[7:0])
    );
    
    acc u_acc_row6_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][1]),
        .acc_data(c1_data[6][15:8]),
        .load_vld(sys_arr_row6_load_vld[1]),
        .load_data(sys_arr_row6_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row6_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row6_data[15:8])
    );
    
    acc u_acc_row6_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][2]),
        .acc_data(c1_data[6][23:16]),
        .load_vld(sys_arr_row6_load_vld[2]),
        .load_data(sys_arr_row6_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row6_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row6_data[23:16])
    );
    
    acc u_acc_row6_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][3]),
        .acc_data(c1_data[6][31:24]),
        .load_vld(sys_arr_row6_load_vld[3]),
        .load_data(sys_arr_row6_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row6_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row6_data[31:24])
    );
    
    acc u_acc_row6_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][4]),
        .acc_data(c1_data[6][39:32]),
        .load_vld(sys_arr_row6_load_vld[4]),
        .load_data(sys_arr_row6_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row6_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row6_data[39:32])
    );
    
    acc u_acc_row6_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][5]),
        .acc_data(c1_data[6][47:40]),
        .load_vld(sys_arr_row6_load_vld[5]),
        .load_data(sys_arr_row6_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row6_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row6_data[47:40])
    );
    
    acc u_acc_row6_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][6]),
        .acc_data(c1_data[6][55:48]),
        .load_vld(sys_arr_row6_load_vld[6]),
        .load_data(sys_arr_row6_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row6_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row6_data[55:48])
    );
    
    acc u_acc_row6_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][7]),
        .acc_data(c1_data[6][63:56]),
        .load_vld(sys_arr_row6_load_vld[7]),
        .load_data(sys_arr_row6_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row6_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row6_data[63:56])
    );
    
    acc u_acc_row6_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][8]),
        .acc_data(c1_data[6][71:64]),
        .load_vld(sys_arr_row6_load_vld[8]),
        .load_data(sys_arr_row6_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row6_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row6_data[71:64])
    );
    
    acc u_acc_row6_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][9]),
        .acc_data(c1_data[6][79:72]),
        .load_vld(sys_arr_row6_load_vld[9]),
        .load_data(sys_arr_row6_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row6_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row6_data[79:72])
    );
    
    acc u_acc_row6_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][10]),
        .acc_data(c1_data[6][87:80]),
        .load_vld(sys_arr_row6_load_vld[10]),
        .load_data(sys_arr_row6_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row6_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row6_data[87:80])
    );
    
    acc u_acc_row6_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][11]),
        .acc_data(c1_data[6][95:88]),
        .load_vld(sys_arr_row6_load_vld[11]),
        .load_data(sys_arr_row6_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row6_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row6_data[95:88])
    );
    
    acc u_acc_row6_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][12]),
        .acc_data(c1_data[6][103:96]),
        .load_vld(sys_arr_row6_load_vld[12]),
        .load_data(sys_arr_row6_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row6_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row6_data[103:96])
    );
    
    acc u_acc_row6_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][13]),
        .acc_data(c1_data[6][111:104]),
        .load_vld(sys_arr_row6_load_vld[13]),
        .load_data(sys_arr_row6_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row6_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row6_data[111:104])
    );
    
    acc u_acc_row6_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][14]),
        .acc_data(c1_data[6][119:112]),
        .load_vld(sys_arr_row6_load_vld[14]),
        .load_data(sys_arr_row6_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row6_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row6_data[119:112])
    );
    
    acc u_acc_row6_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[6][15]),
        .acc_data(c1_data[6][127:120]),
        .load_vld(sys_arr_row6_load_vld[15]),
        .load_data(sys_arr_row6_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row6_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row6_data[127:120])
    );
    
    acc u_acc_row7_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][0]),
        .acc_data(c1_data[7][7:0]),
        .load_vld(sys_arr_row7_load_vld[0]),
        .load_data(sys_arr_row7_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row7_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row7_data[7:0])
    );
    
    acc u_acc_row7_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][1]),
        .acc_data(c1_data[7][15:8]),
        .load_vld(sys_arr_row7_load_vld[1]),
        .load_data(sys_arr_row7_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row7_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row7_data[15:8])
    );
    
    acc u_acc_row7_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][2]),
        .acc_data(c1_data[7][23:16]),
        .load_vld(sys_arr_row7_load_vld[2]),
        .load_data(sys_arr_row7_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row7_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row7_data[23:16])
    );
    
    acc u_acc_row7_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][3]),
        .acc_data(c1_data[7][31:24]),
        .load_vld(sys_arr_row7_load_vld[3]),
        .load_data(sys_arr_row7_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row7_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row7_data[31:24])
    );
    
    acc u_acc_row7_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][4]),
        .acc_data(c1_data[7][39:32]),
        .load_vld(sys_arr_row7_load_vld[4]),
        .load_data(sys_arr_row7_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row7_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row7_data[39:32])
    );
    
    acc u_acc_row7_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][5]),
        .acc_data(c1_data[7][47:40]),
        .load_vld(sys_arr_row7_load_vld[5]),
        .load_data(sys_arr_row7_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row7_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row7_data[47:40])
    );
    
    acc u_acc_row7_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][6]),
        .acc_data(c1_data[7][55:48]),
        .load_vld(sys_arr_row7_load_vld[6]),
        .load_data(sys_arr_row7_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row7_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row7_data[55:48])
    );
    
    acc u_acc_row7_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][7]),
        .acc_data(c1_data[7][63:56]),
        .load_vld(sys_arr_row7_load_vld[7]),
        .load_data(sys_arr_row7_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row7_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row7_data[63:56])
    );
    
    acc u_acc_row7_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][8]),
        .acc_data(c1_data[7][71:64]),
        .load_vld(sys_arr_row7_load_vld[8]),
        .load_data(sys_arr_row7_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row7_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row7_data[71:64])
    );
    
    acc u_acc_row7_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][9]),
        .acc_data(c1_data[7][79:72]),
        .load_vld(sys_arr_row7_load_vld[9]),
        .load_data(sys_arr_row7_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row7_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row7_data[79:72])
    );
    
    acc u_acc_row7_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][10]),
        .acc_data(c1_data[7][87:80]),
        .load_vld(sys_arr_row7_load_vld[10]),
        .load_data(sys_arr_row7_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row7_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row7_data[87:80])
    );
    
    acc u_acc_row7_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][11]),
        .acc_data(c1_data[7][95:88]),
        .load_vld(sys_arr_row7_load_vld[11]),
        .load_data(sys_arr_row7_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row7_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row7_data[95:88])
    );
    
    acc u_acc_row7_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][12]),
        .acc_data(c1_data[7][103:96]),
        .load_vld(sys_arr_row7_load_vld[12]),
        .load_data(sys_arr_row7_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row7_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row7_data[103:96])
    );
    
    acc u_acc_row7_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][13]),
        .acc_data(c1_data[7][111:104]),
        .load_vld(sys_arr_row7_load_vld[13]),
        .load_data(sys_arr_row7_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row7_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row7_data[111:104])
    );
    
    acc u_acc_row7_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][14]),
        .acc_data(c1_data[7][119:112]),
        .load_vld(sys_arr_row7_load_vld[14]),
        .load_data(sys_arr_row7_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row7_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row7_data[119:112])
    );
    
    acc u_acc_row7_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[7][15]),
        .acc_data(c1_data[7][127:120]),
        .load_vld(sys_arr_row7_load_vld[15]),
        .load_data(sys_arr_row7_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row7_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row7_data[127:120])
    );
    
    acc u_acc_row8_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][0]),
        .acc_data(c1_data[8][7:0]),
        .load_vld(sys_arr_row8_load_vld[0]),
        .load_data(sys_arr_row8_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row8_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row8_data[7:0])
    );
    
    acc u_acc_row8_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][1]),
        .acc_data(c1_data[8][15:8]),
        .load_vld(sys_arr_row8_load_vld[1]),
        .load_data(sys_arr_row8_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row8_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row8_data[15:8])
    );
    
    acc u_acc_row8_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][2]),
        .acc_data(c1_data[8][23:16]),
        .load_vld(sys_arr_row8_load_vld[2]),
        .load_data(sys_arr_row8_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row8_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row8_data[23:16])
    );
    
    acc u_acc_row8_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][3]),
        .acc_data(c1_data[8][31:24]),
        .load_vld(sys_arr_row8_load_vld[3]),
        .load_data(sys_arr_row8_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row8_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row8_data[31:24])
    );
    
    acc u_acc_row8_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][4]),
        .acc_data(c1_data[8][39:32]),
        .load_vld(sys_arr_row8_load_vld[4]),
        .load_data(sys_arr_row8_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row8_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row8_data[39:32])
    );
    
    acc u_acc_row8_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][5]),
        .acc_data(c1_data[8][47:40]),
        .load_vld(sys_arr_row8_load_vld[5]),
        .load_data(sys_arr_row8_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row8_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row8_data[47:40])
    );
    
    acc u_acc_row8_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][6]),
        .acc_data(c1_data[8][55:48]),
        .load_vld(sys_arr_row8_load_vld[6]),
        .load_data(sys_arr_row8_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row8_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row8_data[55:48])
    );
    
    acc u_acc_row8_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][7]),
        .acc_data(c1_data[8][63:56]),
        .load_vld(sys_arr_row8_load_vld[7]),
        .load_data(sys_arr_row8_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row8_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row8_data[63:56])
    );
    
    acc u_acc_row8_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][8]),
        .acc_data(c1_data[8][71:64]),
        .load_vld(sys_arr_row8_load_vld[8]),
        .load_data(sys_arr_row8_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row8_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row8_data[71:64])
    );
    
    acc u_acc_row8_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][9]),
        .acc_data(c1_data[8][79:72]),
        .load_vld(sys_arr_row8_load_vld[9]),
        .load_data(sys_arr_row8_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row8_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row8_data[79:72])
    );
    
    acc u_acc_row8_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][10]),
        .acc_data(c1_data[8][87:80]),
        .load_vld(sys_arr_row8_load_vld[10]),
        .load_data(sys_arr_row8_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row8_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row8_data[87:80])
    );
    
    acc u_acc_row8_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][11]),
        .acc_data(c1_data[8][95:88]),
        .load_vld(sys_arr_row8_load_vld[11]),
        .load_data(sys_arr_row8_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row8_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row8_data[95:88])
    );
    
    acc u_acc_row8_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][12]),
        .acc_data(c1_data[8][103:96]),
        .load_vld(sys_arr_row8_load_vld[12]),
        .load_data(sys_arr_row8_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row8_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row8_data[103:96])
    );
    
    acc u_acc_row8_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][13]),
        .acc_data(c1_data[8][111:104]),
        .load_vld(sys_arr_row8_load_vld[13]),
        .load_data(sys_arr_row8_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row8_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row8_data[111:104])
    );
    
    acc u_acc_row8_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][14]),
        .acc_data(c1_data[8][119:112]),
        .load_vld(sys_arr_row8_load_vld[14]),
        .load_data(sys_arr_row8_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row8_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row8_data[119:112])
    );
    
    acc u_acc_row8_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[8][15]),
        .acc_data(c1_data[8][127:120]),
        .load_vld(sys_arr_row8_load_vld[15]),
        .load_data(sys_arr_row8_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row8_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row8_data[127:120])
    );
    
    acc u_acc_row9_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][0]),
        .acc_data(c1_data[9][7:0]),
        .load_vld(sys_arr_row9_load_vld[0]),
        .load_data(sys_arr_row9_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row9_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row9_data[7:0])
    );
    
    acc u_acc_row9_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][1]),
        .acc_data(c1_data[9][15:8]),
        .load_vld(sys_arr_row9_load_vld[1]),
        .load_data(sys_arr_row9_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row9_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row9_data[15:8])
    );
    
    acc u_acc_row9_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][2]),
        .acc_data(c1_data[9][23:16]),
        .load_vld(sys_arr_row9_load_vld[2]),
        .load_data(sys_arr_row9_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row9_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row9_data[23:16])
    );
    
    acc u_acc_row9_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][3]),
        .acc_data(c1_data[9][31:24]),
        .load_vld(sys_arr_row9_load_vld[3]),
        .load_data(sys_arr_row9_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row9_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row9_data[31:24])
    );
    
    acc u_acc_row9_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][4]),
        .acc_data(c1_data[9][39:32]),
        .load_vld(sys_arr_row9_load_vld[4]),
        .load_data(sys_arr_row9_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row9_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row9_data[39:32])
    );
    
    acc u_acc_row9_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][5]),
        .acc_data(c1_data[9][47:40]),
        .load_vld(sys_arr_row9_load_vld[5]),
        .load_data(sys_arr_row9_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row9_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row9_data[47:40])
    );
    
    acc u_acc_row9_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][6]),
        .acc_data(c1_data[9][55:48]),
        .load_vld(sys_arr_row9_load_vld[6]),
        .load_data(sys_arr_row9_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row9_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row9_data[55:48])
    );
    
    acc u_acc_row9_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][7]),
        .acc_data(c1_data[9][63:56]),
        .load_vld(sys_arr_row9_load_vld[7]),
        .load_data(sys_arr_row9_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row9_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row9_data[63:56])
    );
    
    acc u_acc_row9_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][8]),
        .acc_data(c1_data[9][71:64]),
        .load_vld(sys_arr_row9_load_vld[8]),
        .load_data(sys_arr_row9_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row9_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row9_data[71:64])
    );
    
    acc u_acc_row9_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][9]),
        .acc_data(c1_data[9][79:72]),
        .load_vld(sys_arr_row9_load_vld[9]),
        .load_data(sys_arr_row9_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row9_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row9_data[79:72])
    );
    
    acc u_acc_row9_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][10]),
        .acc_data(c1_data[9][87:80]),
        .load_vld(sys_arr_row9_load_vld[10]),
        .load_data(sys_arr_row9_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row9_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row9_data[87:80])
    );
    
    acc u_acc_row9_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][11]),
        .acc_data(c1_data[9][95:88]),
        .load_vld(sys_arr_row9_load_vld[11]),
        .load_data(sys_arr_row9_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row9_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row9_data[95:88])
    );
    
    acc u_acc_row9_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][12]),
        .acc_data(c1_data[9][103:96]),
        .load_vld(sys_arr_row9_load_vld[12]),
        .load_data(sys_arr_row9_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row9_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row9_data[103:96])
    );
    
    acc u_acc_row9_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][13]),
        .acc_data(c1_data[9][111:104]),
        .load_vld(sys_arr_row9_load_vld[13]),
        .load_data(sys_arr_row9_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row9_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row9_data[111:104])
    );
    
    acc u_acc_row9_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][14]),
        .acc_data(c1_data[9][119:112]),
        .load_vld(sys_arr_row9_load_vld[14]),
        .load_data(sys_arr_row9_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row9_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row9_data[119:112])
    );
    
    acc u_acc_row9_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[9][15]),
        .acc_data(c1_data[9][127:120]),
        .load_vld(sys_arr_row9_load_vld[15]),
        .load_data(sys_arr_row9_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row9_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row9_data[127:120])
    );
    
    acc u_acc_row10_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][0]),
        .acc_data(c1_data[10][7:0]),
        .load_vld(sys_arr_row10_load_vld[0]),
        .load_data(sys_arr_row10_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row10_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row10_data[7:0])
    );
    
    acc u_acc_row10_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][1]),
        .acc_data(c1_data[10][15:8]),
        .load_vld(sys_arr_row10_load_vld[1]),
        .load_data(sys_arr_row10_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row10_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row10_data[15:8])
    );
    
    acc u_acc_row10_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][2]),
        .acc_data(c1_data[10][23:16]),
        .load_vld(sys_arr_row10_load_vld[2]),
        .load_data(sys_arr_row10_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row10_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row10_data[23:16])
    );
    
    acc u_acc_row10_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][3]),
        .acc_data(c1_data[10][31:24]),
        .load_vld(sys_arr_row10_load_vld[3]),
        .load_data(sys_arr_row10_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row10_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row10_data[31:24])
    );
    
    acc u_acc_row10_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][4]),
        .acc_data(c1_data[10][39:32]),
        .load_vld(sys_arr_row10_load_vld[4]),
        .load_data(sys_arr_row10_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row10_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row10_data[39:32])
    );
    
    acc u_acc_row10_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][5]),
        .acc_data(c1_data[10][47:40]),
        .load_vld(sys_arr_row10_load_vld[5]),
        .load_data(sys_arr_row10_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row10_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row10_data[47:40])
    );
    
    acc u_acc_row10_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][6]),
        .acc_data(c1_data[10][55:48]),
        .load_vld(sys_arr_row10_load_vld[6]),
        .load_data(sys_arr_row10_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row10_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row10_data[55:48])
    );
    
    acc u_acc_row10_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][7]),
        .acc_data(c1_data[10][63:56]),
        .load_vld(sys_arr_row10_load_vld[7]),
        .load_data(sys_arr_row10_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row10_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row10_data[63:56])
    );
    
    acc u_acc_row10_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][8]),
        .acc_data(c1_data[10][71:64]),
        .load_vld(sys_arr_row10_load_vld[8]),
        .load_data(sys_arr_row10_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row10_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row10_data[71:64])
    );
    
    acc u_acc_row10_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][9]),
        .acc_data(c1_data[10][79:72]),
        .load_vld(sys_arr_row10_load_vld[9]),
        .load_data(sys_arr_row10_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row10_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row10_data[79:72])
    );
    
    acc u_acc_row10_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][10]),
        .acc_data(c1_data[10][87:80]),
        .load_vld(sys_arr_row10_load_vld[10]),
        .load_data(sys_arr_row10_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row10_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row10_data[87:80])
    );
    
    acc u_acc_row10_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][11]),
        .acc_data(c1_data[10][95:88]),
        .load_vld(sys_arr_row10_load_vld[11]),
        .load_data(sys_arr_row10_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row10_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row10_data[95:88])
    );
    
    acc u_acc_row10_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][12]),
        .acc_data(c1_data[10][103:96]),
        .load_vld(sys_arr_row10_load_vld[12]),
        .load_data(sys_arr_row10_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row10_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row10_data[103:96])
    );
    
    acc u_acc_row10_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][13]),
        .acc_data(c1_data[10][111:104]),
        .load_vld(sys_arr_row10_load_vld[13]),
        .load_data(sys_arr_row10_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row10_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row10_data[111:104])
    );
    
    acc u_acc_row10_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][14]),
        .acc_data(c1_data[10][119:112]),
        .load_vld(sys_arr_row10_load_vld[14]),
        .load_data(sys_arr_row10_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row10_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row10_data[119:112])
    );
    
    acc u_acc_row10_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[10][15]),
        .acc_data(c1_data[10][127:120]),
        .load_vld(sys_arr_row10_load_vld[15]),
        .load_data(sys_arr_row10_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row10_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row10_data[127:120])
    );
    
    acc u_acc_row11_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][0]),
        .acc_data(c1_data[11][7:0]),
        .load_vld(sys_arr_row11_load_vld[0]),
        .load_data(sys_arr_row11_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row11_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row11_data[7:0])
    );
    
    acc u_acc_row11_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][1]),
        .acc_data(c1_data[11][15:8]),
        .load_vld(sys_arr_row11_load_vld[1]),
        .load_data(sys_arr_row11_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row11_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row11_data[15:8])
    );
    
    acc u_acc_row11_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][2]),
        .acc_data(c1_data[11][23:16]),
        .load_vld(sys_arr_row11_load_vld[2]),
        .load_data(sys_arr_row11_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row11_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row11_data[23:16])
    );
    
    acc u_acc_row11_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][3]),
        .acc_data(c1_data[11][31:24]),
        .load_vld(sys_arr_row11_load_vld[3]),
        .load_data(sys_arr_row11_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row11_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row11_data[31:24])
    );
    
    acc u_acc_row11_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][4]),
        .acc_data(c1_data[11][39:32]),
        .load_vld(sys_arr_row11_load_vld[4]),
        .load_data(sys_arr_row11_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row11_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row11_data[39:32])
    );
    
    acc u_acc_row11_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][5]),
        .acc_data(c1_data[11][47:40]),
        .load_vld(sys_arr_row11_load_vld[5]),
        .load_data(sys_arr_row11_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row11_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row11_data[47:40])
    );
    
    acc u_acc_row11_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][6]),
        .acc_data(c1_data[11][55:48]),
        .load_vld(sys_arr_row11_load_vld[6]),
        .load_data(sys_arr_row11_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row11_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row11_data[55:48])
    );
    
    acc u_acc_row11_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][7]),
        .acc_data(c1_data[11][63:56]),
        .load_vld(sys_arr_row11_load_vld[7]),
        .load_data(sys_arr_row11_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row11_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row11_data[63:56])
    );
    
    acc u_acc_row11_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][8]),
        .acc_data(c1_data[11][71:64]),
        .load_vld(sys_arr_row11_load_vld[8]),
        .load_data(sys_arr_row11_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row11_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row11_data[71:64])
    );
    
    acc u_acc_row11_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][9]),
        .acc_data(c1_data[11][79:72]),
        .load_vld(sys_arr_row11_load_vld[9]),
        .load_data(sys_arr_row11_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row11_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row11_data[79:72])
    );
    
    acc u_acc_row11_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][10]),
        .acc_data(c1_data[11][87:80]),
        .load_vld(sys_arr_row11_load_vld[10]),
        .load_data(sys_arr_row11_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row11_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row11_data[87:80])
    );
    
    acc u_acc_row11_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][11]),
        .acc_data(c1_data[11][95:88]),
        .load_vld(sys_arr_row11_load_vld[11]),
        .load_data(sys_arr_row11_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row11_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row11_data[95:88])
    );
    
    acc u_acc_row11_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][12]),
        .acc_data(c1_data[11][103:96]),
        .load_vld(sys_arr_row11_load_vld[12]),
        .load_data(sys_arr_row11_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row11_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row11_data[103:96])
    );
    
    acc u_acc_row11_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][13]),
        .acc_data(c1_data[11][111:104]),
        .load_vld(sys_arr_row11_load_vld[13]),
        .load_data(sys_arr_row11_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row11_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row11_data[111:104])
    );
    
    acc u_acc_row11_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][14]),
        .acc_data(c1_data[11][119:112]),
        .load_vld(sys_arr_row11_load_vld[14]),
        .load_data(sys_arr_row11_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row11_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row11_data[119:112])
    );
    
    acc u_acc_row11_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[11][15]),
        .acc_data(c1_data[11][127:120]),
        .load_vld(sys_arr_row11_load_vld[15]),
        .load_data(sys_arr_row11_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row11_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row11_data[127:120])
    );
    
    acc u_acc_row12_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][0]),
        .acc_data(c1_data[12][7:0]),
        .load_vld(sys_arr_row12_load_vld[0]),
        .load_data(sys_arr_row12_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row12_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row12_data[7:0])
    );
    
    acc u_acc_row12_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][1]),
        .acc_data(c1_data[12][15:8]),
        .load_vld(sys_arr_row12_load_vld[1]),
        .load_data(sys_arr_row12_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row12_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row12_data[15:8])
    );
    
    acc u_acc_row12_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][2]),
        .acc_data(c1_data[12][23:16]),
        .load_vld(sys_arr_row12_load_vld[2]),
        .load_data(sys_arr_row12_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row12_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row12_data[23:16])
    );
    
    acc u_acc_row12_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][3]),
        .acc_data(c1_data[12][31:24]),
        .load_vld(sys_arr_row12_load_vld[3]),
        .load_data(sys_arr_row12_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row12_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row12_data[31:24])
    );
    
    acc u_acc_row12_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][4]),
        .acc_data(c1_data[12][39:32]),
        .load_vld(sys_arr_row12_load_vld[4]),
        .load_data(sys_arr_row12_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row12_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row12_data[39:32])
    );
    
    acc u_acc_row12_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][5]),
        .acc_data(c1_data[12][47:40]),
        .load_vld(sys_arr_row12_load_vld[5]),
        .load_data(sys_arr_row12_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row12_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row12_data[47:40])
    );
    
    acc u_acc_row12_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][6]),
        .acc_data(c1_data[12][55:48]),
        .load_vld(sys_arr_row12_load_vld[6]),
        .load_data(sys_arr_row12_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row12_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row12_data[55:48])
    );
    
    acc u_acc_row12_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][7]),
        .acc_data(c1_data[12][63:56]),
        .load_vld(sys_arr_row12_load_vld[7]),
        .load_data(sys_arr_row12_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row12_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row12_data[63:56])
    );
    
    acc u_acc_row12_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][8]),
        .acc_data(c1_data[12][71:64]),
        .load_vld(sys_arr_row12_load_vld[8]),
        .load_data(sys_arr_row12_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row12_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row12_data[71:64])
    );
    
    acc u_acc_row12_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][9]),
        .acc_data(c1_data[12][79:72]),
        .load_vld(sys_arr_row12_load_vld[9]),
        .load_data(sys_arr_row12_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row12_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row12_data[79:72])
    );
    
    acc u_acc_row12_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][10]),
        .acc_data(c1_data[12][87:80]),
        .load_vld(sys_arr_row12_load_vld[10]),
        .load_data(sys_arr_row12_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row12_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row12_data[87:80])
    );
    
    acc u_acc_row12_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][11]),
        .acc_data(c1_data[12][95:88]),
        .load_vld(sys_arr_row12_load_vld[11]),
        .load_data(sys_arr_row12_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row12_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row12_data[95:88])
    );
    
    acc u_acc_row12_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][12]),
        .acc_data(c1_data[12][103:96]),
        .load_vld(sys_arr_row12_load_vld[12]),
        .load_data(sys_arr_row12_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row12_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row12_data[103:96])
    );
    
    acc u_acc_row12_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][13]),
        .acc_data(c1_data[12][111:104]),
        .load_vld(sys_arr_row12_load_vld[13]),
        .load_data(sys_arr_row12_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row12_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row12_data[111:104])
    );
    
    acc u_acc_row12_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][14]),
        .acc_data(c1_data[12][119:112]),
        .load_vld(sys_arr_row12_load_vld[14]),
        .load_data(sys_arr_row12_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row12_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row12_data[119:112])
    );
    
    acc u_acc_row12_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[12][15]),
        .acc_data(c1_data[12][127:120]),
        .load_vld(sys_arr_row12_load_vld[15]),
        .load_data(sys_arr_row12_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row12_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row12_data[127:120])
    );
    
    acc u_acc_row13_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][0]),
        .acc_data(c1_data[13][7:0]),
        .load_vld(sys_arr_row13_load_vld[0]),
        .load_data(sys_arr_row13_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row13_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row13_data[7:0])
    );
    
    acc u_acc_row13_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][1]),
        .acc_data(c1_data[13][15:8]),
        .load_vld(sys_arr_row13_load_vld[1]),
        .load_data(sys_arr_row13_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row13_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row13_data[15:8])
    );
    
    acc u_acc_row13_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][2]),
        .acc_data(c1_data[13][23:16]),
        .load_vld(sys_arr_row13_load_vld[2]),
        .load_data(sys_arr_row13_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row13_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row13_data[23:16])
    );
    
    acc u_acc_row13_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][3]),
        .acc_data(c1_data[13][31:24]),
        .load_vld(sys_arr_row13_load_vld[3]),
        .load_data(sys_arr_row13_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row13_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row13_data[31:24])
    );
    
    acc u_acc_row13_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][4]),
        .acc_data(c1_data[13][39:32]),
        .load_vld(sys_arr_row13_load_vld[4]),
        .load_data(sys_arr_row13_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row13_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row13_data[39:32])
    );
    
    acc u_acc_row13_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][5]),
        .acc_data(c1_data[13][47:40]),
        .load_vld(sys_arr_row13_load_vld[5]),
        .load_data(sys_arr_row13_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row13_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row13_data[47:40])
    );
    
    acc u_acc_row13_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][6]),
        .acc_data(c1_data[13][55:48]),
        .load_vld(sys_arr_row13_load_vld[6]),
        .load_data(sys_arr_row13_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row13_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row13_data[55:48])
    );
    
    acc u_acc_row13_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][7]),
        .acc_data(c1_data[13][63:56]),
        .load_vld(sys_arr_row13_load_vld[7]),
        .load_data(sys_arr_row13_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row13_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row13_data[63:56])
    );
    
    acc u_acc_row13_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][8]),
        .acc_data(c1_data[13][71:64]),
        .load_vld(sys_arr_row13_load_vld[8]),
        .load_data(sys_arr_row13_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row13_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row13_data[71:64])
    );
    
    acc u_acc_row13_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][9]),
        .acc_data(c1_data[13][79:72]),
        .load_vld(sys_arr_row13_load_vld[9]),
        .load_data(sys_arr_row13_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row13_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row13_data[79:72])
    );
    
    acc u_acc_row13_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][10]),
        .acc_data(c1_data[13][87:80]),
        .load_vld(sys_arr_row13_load_vld[10]),
        .load_data(sys_arr_row13_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row13_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row13_data[87:80])
    );
    
    acc u_acc_row13_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][11]),
        .acc_data(c1_data[13][95:88]),
        .load_vld(sys_arr_row13_load_vld[11]),
        .load_data(sys_arr_row13_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row13_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row13_data[95:88])
    );
    
    acc u_acc_row13_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][12]),
        .acc_data(c1_data[13][103:96]),
        .load_vld(sys_arr_row13_load_vld[12]),
        .load_data(sys_arr_row13_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row13_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row13_data[103:96])
    );
    
    acc u_acc_row13_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][13]),
        .acc_data(c1_data[13][111:104]),
        .load_vld(sys_arr_row13_load_vld[13]),
        .load_data(sys_arr_row13_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row13_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row13_data[111:104])
    );
    
    acc u_acc_row13_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][14]),
        .acc_data(c1_data[13][119:112]),
        .load_vld(sys_arr_row13_load_vld[14]),
        .load_data(sys_arr_row13_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row13_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row13_data[119:112])
    );
    
    acc u_acc_row13_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[13][15]),
        .acc_data(c1_data[13][127:120]),
        .load_vld(sys_arr_row13_load_vld[15]),
        .load_data(sys_arr_row13_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row13_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row13_data[127:120])
    );
    
    acc u_acc_row14_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][0]),
        .acc_data(c1_data[14][7:0]),
        .load_vld(sys_arr_row14_load_vld[0]),
        .load_data(sys_arr_row14_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row14_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row14_data[7:0])
    );
    
    acc u_acc_row14_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][1]),
        .acc_data(c1_data[14][15:8]),
        .load_vld(sys_arr_row14_load_vld[1]),
        .load_data(sys_arr_row14_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row14_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row14_data[15:8])
    );
    
    acc u_acc_row14_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][2]),
        .acc_data(c1_data[14][23:16]),
        .load_vld(sys_arr_row14_load_vld[2]),
        .load_data(sys_arr_row14_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row14_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row14_data[23:16])
    );
    
    acc u_acc_row14_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][3]),
        .acc_data(c1_data[14][31:24]),
        .load_vld(sys_arr_row14_load_vld[3]),
        .load_data(sys_arr_row14_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row14_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row14_data[31:24])
    );
    
    acc u_acc_row14_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][4]),
        .acc_data(c1_data[14][39:32]),
        .load_vld(sys_arr_row14_load_vld[4]),
        .load_data(sys_arr_row14_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row14_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row14_data[39:32])
    );
    
    acc u_acc_row14_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][5]),
        .acc_data(c1_data[14][47:40]),
        .load_vld(sys_arr_row14_load_vld[5]),
        .load_data(sys_arr_row14_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row14_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row14_data[47:40])
    );
    
    acc u_acc_row14_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][6]),
        .acc_data(c1_data[14][55:48]),
        .load_vld(sys_arr_row14_load_vld[6]),
        .load_data(sys_arr_row14_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row14_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row14_data[55:48])
    );
    
    acc u_acc_row14_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][7]),
        .acc_data(c1_data[14][63:56]),
        .load_vld(sys_arr_row14_load_vld[7]),
        .load_data(sys_arr_row14_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row14_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row14_data[63:56])
    );
    
    acc u_acc_row14_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][8]),
        .acc_data(c1_data[14][71:64]),
        .load_vld(sys_arr_row14_load_vld[8]),
        .load_data(sys_arr_row14_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row14_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row14_data[71:64])
    );
    
    acc u_acc_row14_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][9]),
        .acc_data(c1_data[14][79:72]),
        .load_vld(sys_arr_row14_load_vld[9]),
        .load_data(sys_arr_row14_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row14_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row14_data[79:72])
    );
    
    acc u_acc_row14_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][10]),
        .acc_data(c1_data[14][87:80]),
        .load_vld(sys_arr_row14_load_vld[10]),
        .load_data(sys_arr_row14_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row14_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row14_data[87:80])
    );
    
    acc u_acc_row14_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][11]),
        .acc_data(c1_data[14][95:88]),
        .load_vld(sys_arr_row14_load_vld[11]),
        .load_data(sys_arr_row14_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row14_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row14_data[95:88])
    );
    
    acc u_acc_row14_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][12]),
        .acc_data(c1_data[14][103:96]),
        .load_vld(sys_arr_row14_load_vld[12]),
        .load_data(sys_arr_row14_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row14_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row14_data[103:96])
    );
    
    acc u_acc_row14_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][13]),
        .acc_data(c1_data[14][111:104]),
        .load_vld(sys_arr_row14_load_vld[13]),
        .load_data(sys_arr_row14_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row14_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row14_data[111:104])
    );
    
    acc u_acc_row14_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][14]),
        .acc_data(c1_data[14][119:112]),
        .load_vld(sys_arr_row14_load_vld[14]),
        .load_data(sys_arr_row14_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row14_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row14_data[119:112])
    );
    
    acc u_acc_row14_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[14][15]),
        .acc_data(c1_data[14][127:120]),
        .load_vld(sys_arr_row14_load_vld[15]),
        .load_data(sys_arr_row14_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row14_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row14_data[127:120])
    );
    
    acc u_acc_row15_col0 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][0]),
        .acc_data(c1_data[15][7:0]),
        .load_vld(sys_arr_row15_load_vld[0]),
        .load_data(sys_arr_row15_load_data[7:0]);
        .out_data_int16(mxu_lsu_int16_row15_data[15:0]),
        .out_data_int8(mxu_lsu_int8_row15_data[7:0])
    );
    
    acc u_acc_row15_col1 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][1]),
        .acc_data(c1_data[15][15:8]),
        .load_vld(sys_arr_row15_load_vld[1]),
        .load_data(sys_arr_row15_load_data[15:8]);
        .out_data_int16(mxu_lsu_int16_row15_data[31:16]),
        .out_data_int8(mxu_lsu_int8_row15_data[15:8])
    );
    
    acc u_acc_row15_col2 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][2]),
        .acc_data(c1_data[15][23:16]),
        .load_vld(sys_arr_row15_load_vld[2]),
        .load_data(sys_arr_row15_load_data[23:16]);
        .out_data_int16(mxu_lsu_int16_row15_data[47:32]),
        .out_data_int8(mxu_lsu_int8_row15_data[23:16])
    );
    
    acc u_acc_row15_col3 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][3]),
        .acc_data(c1_data[15][31:24]),
        .load_vld(sys_arr_row15_load_vld[3]),
        .load_data(sys_arr_row15_load_data[31:24]);
        .out_data_int16(mxu_lsu_int16_row15_data[63:48]),
        .out_data_int8(mxu_lsu_int8_row15_data[31:24])
    );
    
    acc u_acc_row15_col4 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][4]),
        .acc_data(c1_data[15][39:32]),
        .load_vld(sys_arr_row15_load_vld[4]),
        .load_data(sys_arr_row15_load_data[39:32]);
        .out_data_int16(mxu_lsu_int16_row15_data[79:64]),
        .out_data_int8(mxu_lsu_int8_row15_data[39:32])
    );
    
    acc u_acc_row15_col5 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][5]),
        .acc_data(c1_data[15][47:40]),
        .load_vld(sys_arr_row15_load_vld[5]),
        .load_data(sys_arr_row15_load_data[47:40]);
        .out_data_int16(mxu_lsu_int16_row15_data[95:80]),
        .out_data_int8(mxu_lsu_int8_row15_data[47:40])
    );
    
    acc u_acc_row15_col6 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][6]),
        .acc_data(c1_data[15][55:48]),
        .load_vld(sys_arr_row15_load_vld[6]),
        .load_data(sys_arr_row15_load_data[55:48]);
        .out_data_int16(mxu_lsu_int16_row15_data[111:96]),
        .out_data_int8(mxu_lsu_int8_row15_data[55:48])
    );
    
    acc u_acc_row15_col7 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][7]),
        .acc_data(c1_data[15][63:56]),
        .load_vld(sys_arr_row15_load_vld[7]),
        .load_data(sys_arr_row15_load_data[63:56]);
        .out_data_int16(mxu_lsu_int16_row15_data[127:112]),
        .out_data_int8(mxu_lsu_int8_row15_data[63:56])
    );
    
    acc u_acc_row15_col8 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][8]),
        .acc_data(c1_data[15][71:64]),
        .load_vld(sys_arr_row15_load_vld[8]),
        .load_data(sys_arr_row15_load_data[71:64]);
        .out_data_int16(mxu_lsu_int16_row15_data[143:128]),
        .out_data_int8(mxu_lsu_int8_row15_data[71:64])
    );
    
    acc u_acc_row15_col9 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][9]),
        .acc_data(c1_data[15][79:72]),
        .load_vld(sys_arr_row15_load_vld[9]),
        .load_data(sys_arr_row15_load_data[79:72]);
        .out_data_int16(mxu_lsu_int16_row15_data[159:144]),
        .out_data_int8(mxu_lsu_int8_row15_data[79:72])
    );
    
    acc u_acc_row15_col10 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][10]),
        .acc_data(c1_data[15][87:80]),
        .load_vld(sys_arr_row15_load_vld[10]),
        .load_data(sys_arr_row15_load_data[87:80]);
        .out_data_int16(mxu_lsu_int16_row15_data[175:160]),
        .out_data_int8(mxu_lsu_int8_row15_data[87:80])
    );
    
    acc u_acc_row15_col11 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][11]),
        .acc_data(c1_data[15][95:88]),
        .load_vld(sys_arr_row15_load_vld[11]),
        .load_data(sys_arr_row15_load_data[95:88]);
        .out_data_int16(mxu_lsu_int16_row15_data[191:176]),
        .out_data_int8(mxu_lsu_int8_row15_data[95:88])
    );
    
    acc u_acc_row15_col12 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][12]),
        .acc_data(c1_data[15][103:96]),
        .load_vld(sys_arr_row15_load_vld[12]),
        .load_data(sys_arr_row15_load_data[103:96]);
        .out_data_int16(mxu_lsu_int16_row15_data[207:192]),
        .out_data_int8(mxu_lsu_int8_row15_data[103:96])
    );
    
    acc u_acc_row15_col13 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][13]),
        .acc_data(c1_data[15][111:104]),
        .load_vld(sys_arr_row15_load_vld[13]),
        .load_data(sys_arr_row15_load_data[111:104]);
        .out_data_int16(mxu_lsu_int16_row15_data[223:208]),
        .out_data_int8(mxu_lsu_int8_row15_data[111:104])
    );
    
    acc u_acc_row15_col14 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][14]),
        .acc_data(c1_data[15][119:112]),
        .load_vld(sys_arr_row15_load_vld[14]),
        .load_data(sys_arr_row15_load_data[119:112]);
        .out_data_int16(mxu_lsu_int16_row15_data[239:224]),
        .out_data_int8(mxu_lsu_int8_row15_data[119:112])
    );
    
    acc u_acc_row15_col15 (
        .clk(clk),
        .rst_n(rst_n),
        .acc_clr(acc_clr_qual),
        .acc_vld(c1_vld[15][15]),
        .acc_data(c1_data[15][127:120]),
        .load_vld(sys_arr_row15_load_vld[15]),
        .load_data(sys_arr_row15_load_data[127:120]);
        .out_data_int16(mxu_lsu_int16_row15_data[255:240]),
        .out_data_int8(mxu_lsu_int8_row15_data[127:120])
    );
    

    act_mod u_act_mod(
        .clk(clk),
        .rst_n(rst_n),
        .act_type(lsu_mxu_act_type),
        .act_vld(mxu_act_vld),
        .row0_data(mxu_lsu_int16_row0_data),
        .act_row0_vld(act_vld[0]),
        .act_row0_data(act_data[0]),
        .row1_data(mxu_lsu_int16_row1_data),
        .act_row1_vld(act_vld[1]),
        .act_row1_data(act_data[1]),
        .row2_data(mxu_lsu_int16_row2_data),
        .act_row2_vld(act_vld[2]),
        .act_row2_data(act_data[2]),
        .row3_data(mxu_lsu_int16_row3_data),
        .act_row3_vld(act_vld[3]),
        .act_row3_data(act_data[3]),
        .row4_data(mxu_lsu_int16_row4_data),
        .act_row4_vld(act_vld[4]),
        .act_row4_data(act_data[4]),
        .row5_data(mxu_lsu_int16_row5_data),
        .act_row5_vld(act_vld[5]),
        .act_row5_data(act_data[5]),
        .row6_data(mxu_lsu_int16_row6_data),
        .act_row6_vld(act_vld[6]),
        .act_row6_data(act_data[6]),
        .row7_data(mxu_lsu_int16_row7_data),
        .act_row7_vld(act_vld[7]),
        .act_row7_data(act_data[7]),
        .row8_data(mxu_lsu_int16_row8_data),
        .act_row8_vld(act_vld[8]),
        .act_row8_data(act_data[8]),
        .row9_data(mxu_lsu_int16_row9_data),
        .act_row9_vld(act_vld[9]),
        .act_row9_data(act_data[9]),
        .row10_data(mxu_lsu_int16_row10_data),
        .act_row10_vld(act_vld[10]),
        .act_row10_data(act_data[10]),
        .row11_data(mxu_lsu_int16_row11_data),
        .act_row11_vld(act_vld[11]),
        .act_row11_data(act_data[11]),
        .row12_data(mxu_lsu_int16_row12_data),
        .act_row12_vld(act_vld[12]),
        .act_row12_data(act_data[12]),
        .row13_data(mxu_lsu_int16_row13_data),
        .act_row13_vld(act_vld[13]),
        .act_row13_data(act_data[13]),
        .row14_data(mxu_lsu_int16_row14_data),
        .act_row14_vld(act_vld[14]),
        .act_row14_data(act_data[14]),
        .row15_data(mxu_lsu_int16_row15_data),
        .act_row15_vld(act_vld[15]),
        .act_row15_data(act_data[15]),
        .act_busy(act_busy)
    );


endmodule