class mxu_output_monitor extends uvm_monitor;

    virtual mxu_intf mxu_if;
    int send_cnt;
    uvm_analysis_port #(mxu_tr) ap;

    `uvm_component_utils(mxu_output_monitor)
    function new(string name = "mxu_output_monitor", uvm_component parent = null);
       super.new(name, parent);
    endfunction //new()
    
    extern function void build_phase(uvm_phase phase);
    extern virtual task main_phase(uvm_phase phase);
    
    extern virtual task collect_matrix_out(mxu_tr tr);
    extern virtual function void final_phase(uvm_phase phase);

endclass //mxu_output_monitor extends superClass

function void mxu_output_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual mxu_intf)::get(this, "", "mxu_if", mxu_if))begin
        `uvm_fatal("mxu_output_monitor", "mxu output_monitor fail to get mxu if")
    end
    ap = new("ap", this);
endfunction

task mxu_output_monitor::main_phase(uvm_phase phase);
    mxu_tr tr;

    tr = new("tr");

    while (1) begin 
        this.collect_matrix_out(tr);
        ap.write(tr);
    end

endtask

task mxu_output_monitor::collect_matrix_out(mxu_tr tr);

    while(1)begin
        @(posedge mxu_if.clk);
        if(mxu_if.lsu_mxu_vld & mxu_if.mxu_lsu_rdy) break;
    end

    //tr.clear_result();
    while(1) begin
    @(negedge mxu_if.clk);
    //wait(mxu_if.mxu_lsu_data_rdy & mxu_if.mxu_lsu_rdy) 
        if(mxu_if.mxu_lsu_data_rdy & mxu_if.mxu_lsu_rdy & ~(|{mxu_if.lsu_mxu_iram_vld, mxu_if.lsu_mxu_wram_vld})) begin
            `uvm_info("mxu_output_monitor", "begin collect result", UVM_MEDIUM)
            send_cnt++;
            tr.matrix_result_int16[0][0] = {{16{mxu_if.mxu_lsu_int16_row0_data[15]}},mxu_if.mxu_lsu_int16_row0_data[15:0]};
            tr.matrix_result_int8[0][0] = {{24{mxu_if.mxu_lsu_int8_row0_data[7]}},mxu_if.mxu_lsu_int8_row0_data[7:0]};
            tr.matrix_result_int16[0][1] = {{16{mxu_if.mxu_lsu_int16_row0_data[31]}},mxu_if.mxu_lsu_int16_row0_data[31:16]};
            tr.matrix_result_int8[0][1] = {{24{mxu_if.mxu_lsu_int8_row0_data[15]}},mxu_if.mxu_lsu_int8_row0_data[15:8]};
            tr.matrix_result_int16[0][2] = {{16{mxu_if.mxu_lsu_int16_row0_data[47]}},mxu_if.mxu_lsu_int16_row0_data[47:32]};
            tr.matrix_result_int8[0][2] = {{24{mxu_if.mxu_lsu_int8_row0_data[23]}},mxu_if.mxu_lsu_int8_row0_data[23:16]};
            tr.matrix_result_int16[0][3] = {{16{mxu_if.mxu_lsu_int16_row0_data[63]}},mxu_if.mxu_lsu_int16_row0_data[63:48]};
            tr.matrix_result_int8[0][3] = {{24{mxu_if.mxu_lsu_int8_row0_data[31]}},mxu_if.mxu_lsu_int8_row0_data[31:24]};
            tr.matrix_result_int16[0][4] = {{16{mxu_if.mxu_lsu_int16_row0_data[79]}},mxu_if.mxu_lsu_int16_row0_data[79:64]};
            tr.matrix_result_int8[0][4] = {{24{mxu_if.mxu_lsu_int8_row0_data[39]}},mxu_if.mxu_lsu_int8_row0_data[39:32]};
            tr.matrix_result_int16[0][5] = {{16{mxu_if.mxu_lsu_int16_row0_data[95]}},mxu_if.mxu_lsu_int16_row0_data[95:80]};
            tr.matrix_result_int8[0][5] = {{24{mxu_if.mxu_lsu_int8_row0_data[47]}},mxu_if.mxu_lsu_int8_row0_data[47:40]};
            tr.matrix_result_int16[0][6] = {{16{mxu_if.mxu_lsu_int16_row0_data[111]}},mxu_if.mxu_lsu_int16_row0_data[111:96]};
            tr.matrix_result_int8[0][6] = {{24{mxu_if.mxu_lsu_int8_row0_data[55]}},mxu_if.mxu_lsu_int8_row0_data[55:48]};
            tr.matrix_result_int16[0][7] = {{16{mxu_if.mxu_lsu_int16_row0_data[127]}},mxu_if.mxu_lsu_int16_row0_data[127:112]};
            tr.matrix_result_int8[0][7] = {{24{mxu_if.mxu_lsu_int8_row0_data[63]}},mxu_if.mxu_lsu_int8_row0_data[63:56]};
            tr.matrix_result_int16[0][8] = {{16{mxu_if.mxu_lsu_int16_row0_data[143]}},mxu_if.mxu_lsu_int16_row0_data[143:128]};
            tr.matrix_result_int8[0][8] = {{24{mxu_if.mxu_lsu_int8_row0_data[71]}},mxu_if.mxu_lsu_int8_row0_data[71:64]};
            tr.matrix_result_int16[0][9] = {{16{mxu_if.mxu_lsu_int16_row0_data[159]}},mxu_if.mxu_lsu_int16_row0_data[159:144]};
            tr.matrix_result_int8[0][9] = {{24{mxu_if.mxu_lsu_int8_row0_data[79]}},mxu_if.mxu_lsu_int8_row0_data[79:72]};
            tr.matrix_result_int16[0][10] = {{16{mxu_if.mxu_lsu_int16_row0_data[175]}},mxu_if.mxu_lsu_int16_row0_data[175:160]};
            tr.matrix_result_int8[0][10] = {{24{mxu_if.mxu_lsu_int8_row0_data[87]}},mxu_if.mxu_lsu_int8_row0_data[87:80]};
            tr.matrix_result_int16[0][11] = {{16{mxu_if.mxu_lsu_int16_row0_data[191]}},mxu_if.mxu_lsu_int16_row0_data[191:176]};
            tr.matrix_result_int8[0][11] = {{24{mxu_if.mxu_lsu_int8_row0_data[95]}},mxu_if.mxu_lsu_int8_row0_data[95:88]};
            tr.matrix_result_int16[0][12] = {{16{mxu_if.mxu_lsu_int16_row0_data[207]}},mxu_if.mxu_lsu_int16_row0_data[207:192]};
            tr.matrix_result_int8[0][12] = {{24{mxu_if.mxu_lsu_int8_row0_data[103]}},mxu_if.mxu_lsu_int8_row0_data[103:96]};
            tr.matrix_result_int16[0][13] = {{16{mxu_if.mxu_lsu_int16_row0_data[223]}},mxu_if.mxu_lsu_int16_row0_data[223:208]};
            tr.matrix_result_int8[0][13] = {{24{mxu_if.mxu_lsu_int8_row0_data[111]}},mxu_if.mxu_lsu_int8_row0_data[111:104]};
            tr.matrix_result_int16[0][14] = {{16{mxu_if.mxu_lsu_int16_row0_data[239]}},mxu_if.mxu_lsu_int16_row0_data[239:224]};
            tr.matrix_result_int8[0][14] = {{24{mxu_if.mxu_lsu_int8_row0_data[119]}},mxu_if.mxu_lsu_int8_row0_data[119:112]};
            tr.matrix_result_int16[0][15] = {{16{mxu_if.mxu_lsu_int16_row0_data[255]}},mxu_if.mxu_lsu_int16_row0_data[255:240]};
            tr.matrix_result_int8[0][15] = {{24{mxu_if.mxu_lsu_int8_row0_data[127]}},mxu_if.mxu_lsu_int8_row0_data[127:120]};
            tr.matrix_result_int16[1][0] = {{16{mxu_if.mxu_lsu_int16_row1_data[15]}},mxu_if.mxu_lsu_int16_row1_data[15:0]};
            tr.matrix_result_int8[1][0] = {{24{mxu_if.mxu_lsu_int8_row1_data[7]}},mxu_if.mxu_lsu_int8_row1_data[7:0]};
            tr.matrix_result_int16[1][1] = {{16{mxu_if.mxu_lsu_int16_row1_data[31]}},mxu_if.mxu_lsu_int16_row1_data[31:16]};
            tr.matrix_result_int8[1][1] = {{24{mxu_if.mxu_lsu_int8_row1_data[15]}},mxu_if.mxu_lsu_int8_row1_data[15:8]};
            tr.matrix_result_int16[1][2] = {{16{mxu_if.mxu_lsu_int16_row1_data[47]}},mxu_if.mxu_lsu_int16_row1_data[47:32]};
            tr.matrix_result_int8[1][2] = {{24{mxu_if.mxu_lsu_int8_row1_data[23]}},mxu_if.mxu_lsu_int8_row1_data[23:16]};
            tr.matrix_result_int16[1][3] = {{16{mxu_if.mxu_lsu_int16_row1_data[63]}},mxu_if.mxu_lsu_int16_row1_data[63:48]};
            tr.matrix_result_int8[1][3] = {{24{mxu_if.mxu_lsu_int8_row1_data[31]}},mxu_if.mxu_lsu_int8_row1_data[31:24]};
            tr.matrix_result_int16[1][4] = {{16{mxu_if.mxu_lsu_int16_row1_data[79]}},mxu_if.mxu_lsu_int16_row1_data[79:64]};
            tr.matrix_result_int8[1][4] = {{24{mxu_if.mxu_lsu_int8_row1_data[39]}},mxu_if.mxu_lsu_int8_row1_data[39:32]};
            tr.matrix_result_int16[1][5] = {{16{mxu_if.mxu_lsu_int16_row1_data[95]}},mxu_if.mxu_lsu_int16_row1_data[95:80]};
            tr.matrix_result_int8[1][5] = {{24{mxu_if.mxu_lsu_int8_row1_data[47]}},mxu_if.mxu_lsu_int8_row1_data[47:40]};
            tr.matrix_result_int16[1][6] = {{16{mxu_if.mxu_lsu_int16_row1_data[111]}},mxu_if.mxu_lsu_int16_row1_data[111:96]};
            tr.matrix_result_int8[1][6] = {{24{mxu_if.mxu_lsu_int8_row1_data[55]}},mxu_if.mxu_lsu_int8_row1_data[55:48]};
            tr.matrix_result_int16[1][7] = {{16{mxu_if.mxu_lsu_int16_row1_data[127]}},mxu_if.mxu_lsu_int16_row1_data[127:112]};
            tr.matrix_result_int8[1][7] = {{24{mxu_if.mxu_lsu_int8_row1_data[63]}},mxu_if.mxu_lsu_int8_row1_data[63:56]};
            tr.matrix_result_int16[1][8] = {{16{mxu_if.mxu_lsu_int16_row1_data[143]}},mxu_if.mxu_lsu_int16_row1_data[143:128]};
            tr.matrix_result_int8[1][8] = {{24{mxu_if.mxu_lsu_int8_row1_data[71]}},mxu_if.mxu_lsu_int8_row1_data[71:64]};
            tr.matrix_result_int16[1][9] = {{16{mxu_if.mxu_lsu_int16_row1_data[159]}},mxu_if.mxu_lsu_int16_row1_data[159:144]};
            tr.matrix_result_int8[1][9] = {{24{mxu_if.mxu_lsu_int8_row1_data[79]}},mxu_if.mxu_lsu_int8_row1_data[79:72]};
            tr.matrix_result_int16[1][10] = {{16{mxu_if.mxu_lsu_int16_row1_data[175]}},mxu_if.mxu_lsu_int16_row1_data[175:160]};
            tr.matrix_result_int8[1][10] = {{24{mxu_if.mxu_lsu_int8_row1_data[87]}},mxu_if.mxu_lsu_int8_row1_data[87:80]};
            tr.matrix_result_int16[1][11] = {{16{mxu_if.mxu_lsu_int16_row1_data[191]}},mxu_if.mxu_lsu_int16_row1_data[191:176]};
            tr.matrix_result_int8[1][11] = {{24{mxu_if.mxu_lsu_int8_row1_data[95]}},mxu_if.mxu_lsu_int8_row1_data[95:88]};
            tr.matrix_result_int16[1][12] = {{16{mxu_if.mxu_lsu_int16_row1_data[207]}},mxu_if.mxu_lsu_int16_row1_data[207:192]};
            tr.matrix_result_int8[1][12] = {{24{mxu_if.mxu_lsu_int8_row1_data[103]}},mxu_if.mxu_lsu_int8_row1_data[103:96]};
            tr.matrix_result_int16[1][13] = {{16{mxu_if.mxu_lsu_int16_row1_data[223]}},mxu_if.mxu_lsu_int16_row1_data[223:208]};
            tr.matrix_result_int8[1][13] = {{24{mxu_if.mxu_lsu_int8_row1_data[111]}},mxu_if.mxu_lsu_int8_row1_data[111:104]};
            tr.matrix_result_int16[1][14] = {{16{mxu_if.mxu_lsu_int16_row1_data[239]}},mxu_if.mxu_lsu_int16_row1_data[239:224]};
            tr.matrix_result_int8[1][14] = {{24{mxu_if.mxu_lsu_int8_row1_data[119]}},mxu_if.mxu_lsu_int8_row1_data[119:112]};
            tr.matrix_result_int16[1][15] = {{16{mxu_if.mxu_lsu_int16_row1_data[255]}},mxu_if.mxu_lsu_int16_row1_data[255:240]};
            tr.matrix_result_int8[1][15] = {{24{mxu_if.mxu_lsu_int8_row1_data[127]}},mxu_if.mxu_lsu_int8_row1_data[127:120]};
            tr.matrix_result_int16[2][0] = {{16{mxu_if.mxu_lsu_int16_row2_data[15]}},mxu_if.mxu_lsu_int16_row2_data[15:0]};
            tr.matrix_result_int8[2][0] = {{24{mxu_if.mxu_lsu_int8_row2_data[7]}},mxu_if.mxu_lsu_int8_row2_data[7:0]};
            tr.matrix_result_int16[2][1] = {{16{mxu_if.mxu_lsu_int16_row2_data[31]}},mxu_if.mxu_lsu_int16_row2_data[31:16]};
            tr.matrix_result_int8[2][1] = {{24{mxu_if.mxu_lsu_int8_row2_data[15]}},mxu_if.mxu_lsu_int8_row2_data[15:8]};
            tr.matrix_result_int16[2][2] = {{16{mxu_if.mxu_lsu_int16_row2_data[47]}},mxu_if.mxu_lsu_int16_row2_data[47:32]};
            tr.matrix_result_int8[2][2] = {{24{mxu_if.mxu_lsu_int8_row2_data[23]}},mxu_if.mxu_lsu_int8_row2_data[23:16]};
            tr.matrix_result_int16[2][3] = {{16{mxu_if.mxu_lsu_int16_row2_data[63]}},mxu_if.mxu_lsu_int16_row2_data[63:48]};
            tr.matrix_result_int8[2][3] = {{24{mxu_if.mxu_lsu_int8_row2_data[31]}},mxu_if.mxu_lsu_int8_row2_data[31:24]};
            tr.matrix_result_int16[2][4] = {{16{mxu_if.mxu_lsu_int16_row2_data[79]}},mxu_if.mxu_lsu_int16_row2_data[79:64]};
            tr.matrix_result_int8[2][4] = {{24{mxu_if.mxu_lsu_int8_row2_data[39]}},mxu_if.mxu_lsu_int8_row2_data[39:32]};
            tr.matrix_result_int16[2][5] = {{16{mxu_if.mxu_lsu_int16_row2_data[95]}},mxu_if.mxu_lsu_int16_row2_data[95:80]};
            tr.matrix_result_int8[2][5] = {{24{mxu_if.mxu_lsu_int8_row2_data[47]}},mxu_if.mxu_lsu_int8_row2_data[47:40]};
            tr.matrix_result_int16[2][6] = {{16{mxu_if.mxu_lsu_int16_row2_data[111]}},mxu_if.mxu_lsu_int16_row2_data[111:96]};
            tr.matrix_result_int8[2][6] = {{24{mxu_if.mxu_lsu_int8_row2_data[55]}},mxu_if.mxu_lsu_int8_row2_data[55:48]};
            tr.matrix_result_int16[2][7] = {{16{mxu_if.mxu_lsu_int16_row2_data[127]}},mxu_if.mxu_lsu_int16_row2_data[127:112]};
            tr.matrix_result_int8[2][7] = {{24{mxu_if.mxu_lsu_int8_row2_data[63]}},mxu_if.mxu_lsu_int8_row2_data[63:56]};
            tr.matrix_result_int16[2][8] = {{16{mxu_if.mxu_lsu_int16_row2_data[143]}},mxu_if.mxu_lsu_int16_row2_data[143:128]};
            tr.matrix_result_int8[2][8] = {{24{mxu_if.mxu_lsu_int8_row2_data[71]}},mxu_if.mxu_lsu_int8_row2_data[71:64]};
            tr.matrix_result_int16[2][9] = {{16{mxu_if.mxu_lsu_int16_row2_data[159]}},mxu_if.mxu_lsu_int16_row2_data[159:144]};
            tr.matrix_result_int8[2][9] = {{24{mxu_if.mxu_lsu_int8_row2_data[79]}},mxu_if.mxu_lsu_int8_row2_data[79:72]};
            tr.matrix_result_int16[2][10] = {{16{mxu_if.mxu_lsu_int16_row2_data[175]}},mxu_if.mxu_lsu_int16_row2_data[175:160]};
            tr.matrix_result_int8[2][10] = {{24{mxu_if.mxu_lsu_int8_row2_data[87]}},mxu_if.mxu_lsu_int8_row2_data[87:80]};
            tr.matrix_result_int16[2][11] = {{16{mxu_if.mxu_lsu_int16_row2_data[191]}},mxu_if.mxu_lsu_int16_row2_data[191:176]};
            tr.matrix_result_int8[2][11] = {{24{mxu_if.mxu_lsu_int8_row2_data[95]}},mxu_if.mxu_lsu_int8_row2_data[95:88]};
            tr.matrix_result_int16[2][12] = {{16{mxu_if.mxu_lsu_int16_row2_data[207]}},mxu_if.mxu_lsu_int16_row2_data[207:192]};
            tr.matrix_result_int8[2][12] = {{24{mxu_if.mxu_lsu_int8_row2_data[103]}},mxu_if.mxu_lsu_int8_row2_data[103:96]};
            tr.matrix_result_int16[2][13] = {{16{mxu_if.mxu_lsu_int16_row2_data[223]}},mxu_if.mxu_lsu_int16_row2_data[223:208]};
            tr.matrix_result_int8[2][13] = {{24{mxu_if.mxu_lsu_int8_row2_data[111]}},mxu_if.mxu_lsu_int8_row2_data[111:104]};
            tr.matrix_result_int16[2][14] = {{16{mxu_if.mxu_lsu_int16_row2_data[239]}},mxu_if.mxu_lsu_int16_row2_data[239:224]};
            tr.matrix_result_int8[2][14] = {{24{mxu_if.mxu_lsu_int8_row2_data[119]}},mxu_if.mxu_lsu_int8_row2_data[119:112]};
            tr.matrix_result_int16[2][15] = {{16{mxu_if.mxu_lsu_int16_row2_data[255]}},mxu_if.mxu_lsu_int16_row2_data[255:240]};
            tr.matrix_result_int8[2][15] = {{24{mxu_if.mxu_lsu_int8_row2_data[127]}},mxu_if.mxu_lsu_int8_row2_data[127:120]};
            tr.matrix_result_int16[3][0] = {{16{mxu_if.mxu_lsu_int16_row3_data[15]}},mxu_if.mxu_lsu_int16_row3_data[15:0]};
            tr.matrix_result_int8[3][0] = {{24{mxu_if.mxu_lsu_int8_row3_data[7]}},mxu_if.mxu_lsu_int8_row3_data[7:0]};
            tr.matrix_result_int16[3][1] = {{16{mxu_if.mxu_lsu_int16_row3_data[31]}},mxu_if.mxu_lsu_int16_row3_data[31:16]};
            tr.matrix_result_int8[3][1] = {{24{mxu_if.mxu_lsu_int8_row3_data[15]}},mxu_if.mxu_lsu_int8_row3_data[15:8]};
            tr.matrix_result_int16[3][2] = {{16{mxu_if.mxu_lsu_int16_row3_data[47]}},mxu_if.mxu_lsu_int16_row3_data[47:32]};
            tr.matrix_result_int8[3][2] = {{24{mxu_if.mxu_lsu_int8_row3_data[23]}},mxu_if.mxu_lsu_int8_row3_data[23:16]};
            tr.matrix_result_int16[3][3] = {{16{mxu_if.mxu_lsu_int16_row3_data[63]}},mxu_if.mxu_lsu_int16_row3_data[63:48]};
            tr.matrix_result_int8[3][3] = {{24{mxu_if.mxu_lsu_int8_row3_data[31]}},mxu_if.mxu_lsu_int8_row3_data[31:24]};
            tr.matrix_result_int16[3][4] = {{16{mxu_if.mxu_lsu_int16_row3_data[79]}},mxu_if.mxu_lsu_int16_row3_data[79:64]};
            tr.matrix_result_int8[3][4] = {{24{mxu_if.mxu_lsu_int8_row3_data[39]}},mxu_if.mxu_lsu_int8_row3_data[39:32]};
            tr.matrix_result_int16[3][5] = {{16{mxu_if.mxu_lsu_int16_row3_data[95]}},mxu_if.mxu_lsu_int16_row3_data[95:80]};
            tr.matrix_result_int8[3][5] = {{24{mxu_if.mxu_lsu_int8_row3_data[47]}},mxu_if.mxu_lsu_int8_row3_data[47:40]};
            tr.matrix_result_int16[3][6] = {{16{mxu_if.mxu_lsu_int16_row3_data[111]}},mxu_if.mxu_lsu_int16_row3_data[111:96]};
            tr.matrix_result_int8[3][6] = {{24{mxu_if.mxu_lsu_int8_row3_data[55]}},mxu_if.mxu_lsu_int8_row3_data[55:48]};
            tr.matrix_result_int16[3][7] = {{16{mxu_if.mxu_lsu_int16_row3_data[127]}},mxu_if.mxu_lsu_int16_row3_data[127:112]};
            tr.matrix_result_int8[3][7] = {{24{mxu_if.mxu_lsu_int8_row3_data[63]}},mxu_if.mxu_lsu_int8_row3_data[63:56]};
            tr.matrix_result_int16[3][8] = {{16{mxu_if.mxu_lsu_int16_row3_data[143]}},mxu_if.mxu_lsu_int16_row3_data[143:128]};
            tr.matrix_result_int8[3][8] = {{24{mxu_if.mxu_lsu_int8_row3_data[71]}},mxu_if.mxu_lsu_int8_row3_data[71:64]};
            tr.matrix_result_int16[3][9] = {{16{mxu_if.mxu_lsu_int16_row3_data[159]}},mxu_if.mxu_lsu_int16_row3_data[159:144]};
            tr.matrix_result_int8[3][9] = {{24{mxu_if.mxu_lsu_int8_row3_data[79]}},mxu_if.mxu_lsu_int8_row3_data[79:72]};
            tr.matrix_result_int16[3][10] = {{16{mxu_if.mxu_lsu_int16_row3_data[175]}},mxu_if.mxu_lsu_int16_row3_data[175:160]};
            tr.matrix_result_int8[3][10] = {{24{mxu_if.mxu_lsu_int8_row3_data[87]}},mxu_if.mxu_lsu_int8_row3_data[87:80]};
            tr.matrix_result_int16[3][11] = {{16{mxu_if.mxu_lsu_int16_row3_data[191]}},mxu_if.mxu_lsu_int16_row3_data[191:176]};
            tr.matrix_result_int8[3][11] = {{24{mxu_if.mxu_lsu_int8_row3_data[95]}},mxu_if.mxu_lsu_int8_row3_data[95:88]};
            tr.matrix_result_int16[3][12] = {{16{mxu_if.mxu_lsu_int16_row3_data[207]}},mxu_if.mxu_lsu_int16_row3_data[207:192]};
            tr.matrix_result_int8[3][12] = {{24{mxu_if.mxu_lsu_int8_row3_data[103]}},mxu_if.mxu_lsu_int8_row3_data[103:96]};
            tr.matrix_result_int16[3][13] = {{16{mxu_if.mxu_lsu_int16_row3_data[223]}},mxu_if.mxu_lsu_int16_row3_data[223:208]};
            tr.matrix_result_int8[3][13] = {{24{mxu_if.mxu_lsu_int8_row3_data[111]}},mxu_if.mxu_lsu_int8_row3_data[111:104]};
            tr.matrix_result_int16[3][14] = {{16{mxu_if.mxu_lsu_int16_row3_data[239]}},mxu_if.mxu_lsu_int16_row3_data[239:224]};
            tr.matrix_result_int8[3][14] = {{24{mxu_if.mxu_lsu_int8_row3_data[119]}},mxu_if.mxu_lsu_int8_row3_data[119:112]};
            tr.matrix_result_int16[3][15] = {{16{mxu_if.mxu_lsu_int16_row3_data[255]}},mxu_if.mxu_lsu_int16_row3_data[255:240]};
            tr.matrix_result_int8[3][15] = {{24{mxu_if.mxu_lsu_int8_row3_data[127]}},mxu_if.mxu_lsu_int8_row3_data[127:120]};
            tr.matrix_result_int16[4][0] = {{16{mxu_if.mxu_lsu_int16_row4_data[15]}},mxu_if.mxu_lsu_int16_row4_data[15:0]};
            tr.matrix_result_int8[4][0] = {{24{mxu_if.mxu_lsu_int8_row4_data[7]}},mxu_if.mxu_lsu_int8_row4_data[7:0]};
            tr.matrix_result_int16[4][1] = {{16{mxu_if.mxu_lsu_int16_row4_data[31]}},mxu_if.mxu_lsu_int16_row4_data[31:16]};
            tr.matrix_result_int8[4][1] = {{24{mxu_if.mxu_lsu_int8_row4_data[15]}},mxu_if.mxu_lsu_int8_row4_data[15:8]};
            tr.matrix_result_int16[4][2] = {{16{mxu_if.mxu_lsu_int16_row4_data[47]}},mxu_if.mxu_lsu_int16_row4_data[47:32]};
            tr.matrix_result_int8[4][2] = {{24{mxu_if.mxu_lsu_int8_row4_data[23]}},mxu_if.mxu_lsu_int8_row4_data[23:16]};
            tr.matrix_result_int16[4][3] = {{16{mxu_if.mxu_lsu_int16_row4_data[63]}},mxu_if.mxu_lsu_int16_row4_data[63:48]};
            tr.matrix_result_int8[4][3] = {{24{mxu_if.mxu_lsu_int8_row4_data[31]}},mxu_if.mxu_lsu_int8_row4_data[31:24]};
            tr.matrix_result_int16[4][4] = {{16{mxu_if.mxu_lsu_int16_row4_data[79]}},mxu_if.mxu_lsu_int16_row4_data[79:64]};
            tr.matrix_result_int8[4][4] = {{24{mxu_if.mxu_lsu_int8_row4_data[39]}},mxu_if.mxu_lsu_int8_row4_data[39:32]};
            tr.matrix_result_int16[4][5] = {{16{mxu_if.mxu_lsu_int16_row4_data[95]}},mxu_if.mxu_lsu_int16_row4_data[95:80]};
            tr.matrix_result_int8[4][5] = {{24{mxu_if.mxu_lsu_int8_row4_data[47]}},mxu_if.mxu_lsu_int8_row4_data[47:40]};
            tr.matrix_result_int16[4][6] = {{16{mxu_if.mxu_lsu_int16_row4_data[111]}},mxu_if.mxu_lsu_int16_row4_data[111:96]};
            tr.matrix_result_int8[4][6] = {{24{mxu_if.mxu_lsu_int8_row4_data[55]}},mxu_if.mxu_lsu_int8_row4_data[55:48]};
            tr.matrix_result_int16[4][7] = {{16{mxu_if.mxu_lsu_int16_row4_data[127]}},mxu_if.mxu_lsu_int16_row4_data[127:112]};
            tr.matrix_result_int8[4][7] = {{24{mxu_if.mxu_lsu_int8_row4_data[63]}},mxu_if.mxu_lsu_int8_row4_data[63:56]};
            tr.matrix_result_int16[4][8] = {{16{mxu_if.mxu_lsu_int16_row4_data[143]}},mxu_if.mxu_lsu_int16_row4_data[143:128]};
            tr.matrix_result_int8[4][8] = {{24{mxu_if.mxu_lsu_int8_row4_data[71]}},mxu_if.mxu_lsu_int8_row4_data[71:64]};
            tr.matrix_result_int16[4][9] = {{16{mxu_if.mxu_lsu_int16_row4_data[159]}},mxu_if.mxu_lsu_int16_row4_data[159:144]};
            tr.matrix_result_int8[4][9] = {{24{mxu_if.mxu_lsu_int8_row4_data[79]}},mxu_if.mxu_lsu_int8_row4_data[79:72]};
            tr.matrix_result_int16[4][10] = {{16{mxu_if.mxu_lsu_int16_row4_data[175]}},mxu_if.mxu_lsu_int16_row4_data[175:160]};
            tr.matrix_result_int8[4][10] = {{24{mxu_if.mxu_lsu_int8_row4_data[87]}},mxu_if.mxu_lsu_int8_row4_data[87:80]};
            tr.matrix_result_int16[4][11] = {{16{mxu_if.mxu_lsu_int16_row4_data[191]}},mxu_if.mxu_lsu_int16_row4_data[191:176]};
            tr.matrix_result_int8[4][11] = {{24{mxu_if.mxu_lsu_int8_row4_data[95]}},mxu_if.mxu_lsu_int8_row4_data[95:88]};
            tr.matrix_result_int16[4][12] = {{16{mxu_if.mxu_lsu_int16_row4_data[207]}},mxu_if.mxu_lsu_int16_row4_data[207:192]};
            tr.matrix_result_int8[4][12] = {{24{mxu_if.mxu_lsu_int8_row4_data[103]}},mxu_if.mxu_lsu_int8_row4_data[103:96]};
            tr.matrix_result_int16[4][13] = {{16{mxu_if.mxu_lsu_int16_row4_data[223]}},mxu_if.mxu_lsu_int16_row4_data[223:208]};
            tr.matrix_result_int8[4][13] = {{24{mxu_if.mxu_lsu_int8_row4_data[111]}},mxu_if.mxu_lsu_int8_row4_data[111:104]};
            tr.matrix_result_int16[4][14] = {{16{mxu_if.mxu_lsu_int16_row4_data[239]}},mxu_if.mxu_lsu_int16_row4_data[239:224]};
            tr.matrix_result_int8[4][14] = {{24{mxu_if.mxu_lsu_int8_row4_data[119]}},mxu_if.mxu_lsu_int8_row4_data[119:112]};
            tr.matrix_result_int16[4][15] = {{16{mxu_if.mxu_lsu_int16_row4_data[255]}},mxu_if.mxu_lsu_int16_row4_data[255:240]};
            tr.matrix_result_int8[4][15] = {{24{mxu_if.mxu_lsu_int8_row4_data[127]}},mxu_if.mxu_lsu_int8_row4_data[127:120]};
            tr.matrix_result_int16[5][0] = {{16{mxu_if.mxu_lsu_int16_row5_data[15]}},mxu_if.mxu_lsu_int16_row5_data[15:0]};
            tr.matrix_result_int8[5][0] = {{24{mxu_if.mxu_lsu_int8_row5_data[7]}},mxu_if.mxu_lsu_int8_row5_data[7:0]};
            tr.matrix_result_int16[5][1] = {{16{mxu_if.mxu_lsu_int16_row5_data[31]}},mxu_if.mxu_lsu_int16_row5_data[31:16]};
            tr.matrix_result_int8[5][1] = {{24{mxu_if.mxu_lsu_int8_row5_data[15]}},mxu_if.mxu_lsu_int8_row5_data[15:8]};
            tr.matrix_result_int16[5][2] = {{16{mxu_if.mxu_lsu_int16_row5_data[47]}},mxu_if.mxu_lsu_int16_row5_data[47:32]};
            tr.matrix_result_int8[5][2] = {{24{mxu_if.mxu_lsu_int8_row5_data[23]}},mxu_if.mxu_lsu_int8_row5_data[23:16]};
            tr.matrix_result_int16[5][3] = {{16{mxu_if.mxu_lsu_int16_row5_data[63]}},mxu_if.mxu_lsu_int16_row5_data[63:48]};
            tr.matrix_result_int8[5][3] = {{24{mxu_if.mxu_lsu_int8_row5_data[31]}},mxu_if.mxu_lsu_int8_row5_data[31:24]};
            tr.matrix_result_int16[5][4] = {{16{mxu_if.mxu_lsu_int16_row5_data[79]}},mxu_if.mxu_lsu_int16_row5_data[79:64]};
            tr.matrix_result_int8[5][4] = {{24{mxu_if.mxu_lsu_int8_row5_data[39]}},mxu_if.mxu_lsu_int8_row5_data[39:32]};
            tr.matrix_result_int16[5][5] = {{16{mxu_if.mxu_lsu_int16_row5_data[95]}},mxu_if.mxu_lsu_int16_row5_data[95:80]};
            tr.matrix_result_int8[5][5] = {{24{mxu_if.mxu_lsu_int8_row5_data[47]}},mxu_if.mxu_lsu_int8_row5_data[47:40]};
            tr.matrix_result_int16[5][6] = {{16{mxu_if.mxu_lsu_int16_row5_data[111]}},mxu_if.mxu_lsu_int16_row5_data[111:96]};
            tr.matrix_result_int8[5][6] = {{24{mxu_if.mxu_lsu_int8_row5_data[55]}},mxu_if.mxu_lsu_int8_row5_data[55:48]};
            tr.matrix_result_int16[5][7] = {{16{mxu_if.mxu_lsu_int16_row5_data[127]}},mxu_if.mxu_lsu_int16_row5_data[127:112]};
            tr.matrix_result_int8[5][7] = {{24{mxu_if.mxu_lsu_int8_row5_data[63]}},mxu_if.mxu_lsu_int8_row5_data[63:56]};
            tr.matrix_result_int16[5][8] = {{16{mxu_if.mxu_lsu_int16_row5_data[143]}},mxu_if.mxu_lsu_int16_row5_data[143:128]};
            tr.matrix_result_int8[5][8] = {{24{mxu_if.mxu_lsu_int8_row5_data[71]}},mxu_if.mxu_lsu_int8_row5_data[71:64]};
            tr.matrix_result_int16[5][9] = {{16{mxu_if.mxu_lsu_int16_row5_data[159]}},mxu_if.mxu_lsu_int16_row5_data[159:144]};
            tr.matrix_result_int8[5][9] = {{24{mxu_if.mxu_lsu_int8_row5_data[79]}},mxu_if.mxu_lsu_int8_row5_data[79:72]};
            tr.matrix_result_int16[5][10] = {{16{mxu_if.mxu_lsu_int16_row5_data[175]}},mxu_if.mxu_lsu_int16_row5_data[175:160]};
            tr.matrix_result_int8[5][10] = {{24{mxu_if.mxu_lsu_int8_row5_data[87]}},mxu_if.mxu_lsu_int8_row5_data[87:80]};
            tr.matrix_result_int16[5][11] = {{16{mxu_if.mxu_lsu_int16_row5_data[191]}},mxu_if.mxu_lsu_int16_row5_data[191:176]};
            tr.matrix_result_int8[5][11] = {{24{mxu_if.mxu_lsu_int8_row5_data[95]}},mxu_if.mxu_lsu_int8_row5_data[95:88]};
            tr.matrix_result_int16[5][12] = {{16{mxu_if.mxu_lsu_int16_row5_data[207]}},mxu_if.mxu_lsu_int16_row5_data[207:192]};
            tr.matrix_result_int8[5][12] = {{24{mxu_if.mxu_lsu_int8_row5_data[103]}},mxu_if.mxu_lsu_int8_row5_data[103:96]};
            tr.matrix_result_int16[5][13] = {{16{mxu_if.mxu_lsu_int16_row5_data[223]}},mxu_if.mxu_lsu_int16_row5_data[223:208]};
            tr.matrix_result_int8[5][13] = {{24{mxu_if.mxu_lsu_int8_row5_data[111]}},mxu_if.mxu_lsu_int8_row5_data[111:104]};
            tr.matrix_result_int16[5][14] = {{16{mxu_if.mxu_lsu_int16_row5_data[239]}},mxu_if.mxu_lsu_int16_row5_data[239:224]};
            tr.matrix_result_int8[5][14] = {{24{mxu_if.mxu_lsu_int8_row5_data[119]}},mxu_if.mxu_lsu_int8_row5_data[119:112]};
            tr.matrix_result_int16[5][15] = {{16{mxu_if.mxu_lsu_int16_row5_data[255]}},mxu_if.mxu_lsu_int16_row5_data[255:240]};
            tr.matrix_result_int8[5][15] = {{24{mxu_if.mxu_lsu_int8_row5_data[127]}},mxu_if.mxu_lsu_int8_row5_data[127:120]};
            tr.matrix_result_int16[6][0] = {{16{mxu_if.mxu_lsu_int16_row6_data[15]}},mxu_if.mxu_lsu_int16_row6_data[15:0]};
            tr.matrix_result_int8[6][0] = {{24{mxu_if.mxu_lsu_int8_row6_data[7]}},mxu_if.mxu_lsu_int8_row6_data[7:0]};
            tr.matrix_result_int16[6][1] = {{16{mxu_if.mxu_lsu_int16_row6_data[31]}},mxu_if.mxu_lsu_int16_row6_data[31:16]};
            tr.matrix_result_int8[6][1] = {{24{mxu_if.mxu_lsu_int8_row6_data[15]}},mxu_if.mxu_lsu_int8_row6_data[15:8]};
            tr.matrix_result_int16[6][2] = {{16{mxu_if.mxu_lsu_int16_row6_data[47]}},mxu_if.mxu_lsu_int16_row6_data[47:32]};
            tr.matrix_result_int8[6][2] = {{24{mxu_if.mxu_lsu_int8_row6_data[23]}},mxu_if.mxu_lsu_int8_row6_data[23:16]};
            tr.matrix_result_int16[6][3] = {{16{mxu_if.mxu_lsu_int16_row6_data[63]}},mxu_if.mxu_lsu_int16_row6_data[63:48]};
            tr.matrix_result_int8[6][3] = {{24{mxu_if.mxu_lsu_int8_row6_data[31]}},mxu_if.mxu_lsu_int8_row6_data[31:24]};
            tr.matrix_result_int16[6][4] = {{16{mxu_if.mxu_lsu_int16_row6_data[79]}},mxu_if.mxu_lsu_int16_row6_data[79:64]};
            tr.matrix_result_int8[6][4] = {{24{mxu_if.mxu_lsu_int8_row6_data[39]}},mxu_if.mxu_lsu_int8_row6_data[39:32]};
            tr.matrix_result_int16[6][5] = {{16{mxu_if.mxu_lsu_int16_row6_data[95]}},mxu_if.mxu_lsu_int16_row6_data[95:80]};
            tr.matrix_result_int8[6][5] = {{24{mxu_if.mxu_lsu_int8_row6_data[47]}},mxu_if.mxu_lsu_int8_row6_data[47:40]};
            tr.matrix_result_int16[6][6] = {{16{mxu_if.mxu_lsu_int16_row6_data[111]}},mxu_if.mxu_lsu_int16_row6_data[111:96]};
            tr.matrix_result_int8[6][6] = {{24{mxu_if.mxu_lsu_int8_row6_data[55]}},mxu_if.mxu_lsu_int8_row6_data[55:48]};
            tr.matrix_result_int16[6][7] = {{16{mxu_if.mxu_lsu_int16_row6_data[127]}},mxu_if.mxu_lsu_int16_row6_data[127:112]};
            tr.matrix_result_int8[6][7] = {{24{mxu_if.mxu_lsu_int8_row6_data[63]}},mxu_if.mxu_lsu_int8_row6_data[63:56]};
            tr.matrix_result_int16[6][8] = {{16{mxu_if.mxu_lsu_int16_row6_data[143]}},mxu_if.mxu_lsu_int16_row6_data[143:128]};
            tr.matrix_result_int8[6][8] = {{24{mxu_if.mxu_lsu_int8_row6_data[71]}},mxu_if.mxu_lsu_int8_row6_data[71:64]};
            tr.matrix_result_int16[6][9] = {{16{mxu_if.mxu_lsu_int16_row6_data[159]}},mxu_if.mxu_lsu_int16_row6_data[159:144]};
            tr.matrix_result_int8[6][9] = {{24{mxu_if.mxu_lsu_int8_row6_data[79]}},mxu_if.mxu_lsu_int8_row6_data[79:72]};
            tr.matrix_result_int16[6][10] = {{16{mxu_if.mxu_lsu_int16_row6_data[175]}},mxu_if.mxu_lsu_int16_row6_data[175:160]};
            tr.matrix_result_int8[6][10] = {{24{mxu_if.mxu_lsu_int8_row6_data[87]}},mxu_if.mxu_lsu_int8_row6_data[87:80]};
            tr.matrix_result_int16[6][11] = {{16{mxu_if.mxu_lsu_int16_row6_data[191]}},mxu_if.mxu_lsu_int16_row6_data[191:176]};
            tr.matrix_result_int8[6][11] = {{24{mxu_if.mxu_lsu_int8_row6_data[95]}},mxu_if.mxu_lsu_int8_row6_data[95:88]};
            tr.matrix_result_int16[6][12] = {{16{mxu_if.mxu_lsu_int16_row6_data[207]}},mxu_if.mxu_lsu_int16_row6_data[207:192]};
            tr.matrix_result_int8[6][12] = {{24{mxu_if.mxu_lsu_int8_row6_data[103]}},mxu_if.mxu_lsu_int8_row6_data[103:96]};
            tr.matrix_result_int16[6][13] = {{16{mxu_if.mxu_lsu_int16_row6_data[223]}},mxu_if.mxu_lsu_int16_row6_data[223:208]};
            tr.matrix_result_int8[6][13] = {{24{mxu_if.mxu_lsu_int8_row6_data[111]}},mxu_if.mxu_lsu_int8_row6_data[111:104]};
            tr.matrix_result_int16[6][14] = {{16{mxu_if.mxu_lsu_int16_row6_data[239]}},mxu_if.mxu_lsu_int16_row6_data[239:224]};
            tr.matrix_result_int8[6][14] = {{24{mxu_if.mxu_lsu_int8_row6_data[119]}},mxu_if.mxu_lsu_int8_row6_data[119:112]};
            tr.matrix_result_int16[6][15] = {{16{mxu_if.mxu_lsu_int16_row6_data[255]}},mxu_if.mxu_lsu_int16_row6_data[255:240]};
            tr.matrix_result_int8[6][15] = {{24{mxu_if.mxu_lsu_int8_row6_data[127]}},mxu_if.mxu_lsu_int8_row6_data[127:120]};
            tr.matrix_result_int16[7][0] = {{16{mxu_if.mxu_lsu_int16_row7_data[15]}},mxu_if.mxu_lsu_int16_row7_data[15:0]};
            tr.matrix_result_int8[7][0] = {{24{mxu_if.mxu_lsu_int8_row7_data[7]}},mxu_if.mxu_lsu_int8_row7_data[7:0]};
            tr.matrix_result_int16[7][1] = {{16{mxu_if.mxu_lsu_int16_row7_data[31]}},mxu_if.mxu_lsu_int16_row7_data[31:16]};
            tr.matrix_result_int8[7][1] = {{24{mxu_if.mxu_lsu_int8_row7_data[15]}},mxu_if.mxu_lsu_int8_row7_data[15:8]};
            tr.matrix_result_int16[7][2] = {{16{mxu_if.mxu_lsu_int16_row7_data[47]}},mxu_if.mxu_lsu_int16_row7_data[47:32]};
            tr.matrix_result_int8[7][2] = {{24{mxu_if.mxu_lsu_int8_row7_data[23]}},mxu_if.mxu_lsu_int8_row7_data[23:16]};
            tr.matrix_result_int16[7][3] = {{16{mxu_if.mxu_lsu_int16_row7_data[63]}},mxu_if.mxu_lsu_int16_row7_data[63:48]};
            tr.matrix_result_int8[7][3] = {{24{mxu_if.mxu_lsu_int8_row7_data[31]}},mxu_if.mxu_lsu_int8_row7_data[31:24]};
            tr.matrix_result_int16[7][4] = {{16{mxu_if.mxu_lsu_int16_row7_data[79]}},mxu_if.mxu_lsu_int16_row7_data[79:64]};
            tr.matrix_result_int8[7][4] = {{24{mxu_if.mxu_lsu_int8_row7_data[39]}},mxu_if.mxu_lsu_int8_row7_data[39:32]};
            tr.matrix_result_int16[7][5] = {{16{mxu_if.mxu_lsu_int16_row7_data[95]}},mxu_if.mxu_lsu_int16_row7_data[95:80]};
            tr.matrix_result_int8[7][5] = {{24{mxu_if.mxu_lsu_int8_row7_data[47]}},mxu_if.mxu_lsu_int8_row7_data[47:40]};
            tr.matrix_result_int16[7][6] = {{16{mxu_if.mxu_lsu_int16_row7_data[111]}},mxu_if.mxu_lsu_int16_row7_data[111:96]};
            tr.matrix_result_int8[7][6] = {{24{mxu_if.mxu_lsu_int8_row7_data[55]}},mxu_if.mxu_lsu_int8_row7_data[55:48]};
            tr.matrix_result_int16[7][7] = {{16{mxu_if.mxu_lsu_int16_row7_data[127]}},mxu_if.mxu_lsu_int16_row7_data[127:112]};
            tr.matrix_result_int8[7][7] = {{24{mxu_if.mxu_lsu_int8_row7_data[63]}},mxu_if.mxu_lsu_int8_row7_data[63:56]};
            tr.matrix_result_int16[7][8] = {{16{mxu_if.mxu_lsu_int16_row7_data[143]}},mxu_if.mxu_lsu_int16_row7_data[143:128]};
            tr.matrix_result_int8[7][8] = {{24{mxu_if.mxu_lsu_int8_row7_data[71]}},mxu_if.mxu_lsu_int8_row7_data[71:64]};
            tr.matrix_result_int16[7][9] = {{16{mxu_if.mxu_lsu_int16_row7_data[159]}},mxu_if.mxu_lsu_int16_row7_data[159:144]};
            tr.matrix_result_int8[7][9] = {{24{mxu_if.mxu_lsu_int8_row7_data[79]}},mxu_if.mxu_lsu_int8_row7_data[79:72]};
            tr.matrix_result_int16[7][10] = {{16{mxu_if.mxu_lsu_int16_row7_data[175]}},mxu_if.mxu_lsu_int16_row7_data[175:160]};
            tr.matrix_result_int8[7][10] = {{24{mxu_if.mxu_lsu_int8_row7_data[87]}},mxu_if.mxu_lsu_int8_row7_data[87:80]};
            tr.matrix_result_int16[7][11] = {{16{mxu_if.mxu_lsu_int16_row7_data[191]}},mxu_if.mxu_lsu_int16_row7_data[191:176]};
            tr.matrix_result_int8[7][11] = {{24{mxu_if.mxu_lsu_int8_row7_data[95]}},mxu_if.mxu_lsu_int8_row7_data[95:88]};
            tr.matrix_result_int16[7][12] = {{16{mxu_if.mxu_lsu_int16_row7_data[207]}},mxu_if.mxu_lsu_int16_row7_data[207:192]};
            tr.matrix_result_int8[7][12] = {{24{mxu_if.mxu_lsu_int8_row7_data[103]}},mxu_if.mxu_lsu_int8_row7_data[103:96]};
            tr.matrix_result_int16[7][13] = {{16{mxu_if.mxu_lsu_int16_row7_data[223]}},mxu_if.mxu_lsu_int16_row7_data[223:208]};
            tr.matrix_result_int8[7][13] = {{24{mxu_if.mxu_lsu_int8_row7_data[111]}},mxu_if.mxu_lsu_int8_row7_data[111:104]};
            tr.matrix_result_int16[7][14] = {{16{mxu_if.mxu_lsu_int16_row7_data[239]}},mxu_if.mxu_lsu_int16_row7_data[239:224]};
            tr.matrix_result_int8[7][14] = {{24{mxu_if.mxu_lsu_int8_row7_data[119]}},mxu_if.mxu_lsu_int8_row7_data[119:112]};
            tr.matrix_result_int16[7][15] = {{16{mxu_if.mxu_lsu_int16_row7_data[255]}},mxu_if.mxu_lsu_int16_row7_data[255:240]};
            tr.matrix_result_int8[7][15] = {{24{mxu_if.mxu_lsu_int8_row7_data[127]}},mxu_if.mxu_lsu_int8_row7_data[127:120]};
            tr.matrix_result_int16[8][0] = {{16{mxu_if.mxu_lsu_int16_row8_data[15]}},mxu_if.mxu_lsu_int16_row8_data[15:0]};
            tr.matrix_result_int8[8][0] = {{24{mxu_if.mxu_lsu_int8_row8_data[7]}},mxu_if.mxu_lsu_int8_row8_data[7:0]};
            tr.matrix_result_int16[8][1] = {{16{mxu_if.mxu_lsu_int16_row8_data[31]}},mxu_if.mxu_lsu_int16_row8_data[31:16]};
            tr.matrix_result_int8[8][1] = {{24{mxu_if.mxu_lsu_int8_row8_data[15]}},mxu_if.mxu_lsu_int8_row8_data[15:8]};
            tr.matrix_result_int16[8][2] = {{16{mxu_if.mxu_lsu_int16_row8_data[47]}},mxu_if.mxu_lsu_int16_row8_data[47:32]};
            tr.matrix_result_int8[8][2] = {{24{mxu_if.mxu_lsu_int8_row8_data[23]}},mxu_if.mxu_lsu_int8_row8_data[23:16]};
            tr.matrix_result_int16[8][3] = {{16{mxu_if.mxu_lsu_int16_row8_data[63]}},mxu_if.mxu_lsu_int16_row8_data[63:48]};
            tr.matrix_result_int8[8][3] = {{24{mxu_if.mxu_lsu_int8_row8_data[31]}},mxu_if.mxu_lsu_int8_row8_data[31:24]};
            tr.matrix_result_int16[8][4] = {{16{mxu_if.mxu_lsu_int16_row8_data[79]}},mxu_if.mxu_lsu_int16_row8_data[79:64]};
            tr.matrix_result_int8[8][4] = {{24{mxu_if.mxu_lsu_int8_row8_data[39]}},mxu_if.mxu_lsu_int8_row8_data[39:32]};
            tr.matrix_result_int16[8][5] = {{16{mxu_if.mxu_lsu_int16_row8_data[95]}},mxu_if.mxu_lsu_int16_row8_data[95:80]};
            tr.matrix_result_int8[8][5] = {{24{mxu_if.mxu_lsu_int8_row8_data[47]}},mxu_if.mxu_lsu_int8_row8_data[47:40]};
            tr.matrix_result_int16[8][6] = {{16{mxu_if.mxu_lsu_int16_row8_data[111]}},mxu_if.mxu_lsu_int16_row8_data[111:96]};
            tr.matrix_result_int8[8][6] = {{24{mxu_if.mxu_lsu_int8_row8_data[55]}},mxu_if.mxu_lsu_int8_row8_data[55:48]};
            tr.matrix_result_int16[8][7] = {{16{mxu_if.mxu_lsu_int16_row8_data[127]}},mxu_if.mxu_lsu_int16_row8_data[127:112]};
            tr.matrix_result_int8[8][7] = {{24{mxu_if.mxu_lsu_int8_row8_data[63]}},mxu_if.mxu_lsu_int8_row8_data[63:56]};
            tr.matrix_result_int16[8][8] = {{16{mxu_if.mxu_lsu_int16_row8_data[143]}},mxu_if.mxu_lsu_int16_row8_data[143:128]};
            tr.matrix_result_int8[8][8] = {{24{mxu_if.mxu_lsu_int8_row8_data[71]}},mxu_if.mxu_lsu_int8_row8_data[71:64]};
            tr.matrix_result_int16[8][9] = {{16{mxu_if.mxu_lsu_int16_row8_data[159]}},mxu_if.mxu_lsu_int16_row8_data[159:144]};
            tr.matrix_result_int8[8][9] = {{24{mxu_if.mxu_lsu_int8_row8_data[79]}},mxu_if.mxu_lsu_int8_row8_data[79:72]};
            tr.matrix_result_int16[8][10] = {{16{mxu_if.mxu_lsu_int16_row8_data[175]}},mxu_if.mxu_lsu_int16_row8_data[175:160]};
            tr.matrix_result_int8[8][10] = {{24{mxu_if.mxu_lsu_int8_row8_data[87]}},mxu_if.mxu_lsu_int8_row8_data[87:80]};
            tr.matrix_result_int16[8][11] = {{16{mxu_if.mxu_lsu_int16_row8_data[191]}},mxu_if.mxu_lsu_int16_row8_data[191:176]};
            tr.matrix_result_int8[8][11] = {{24{mxu_if.mxu_lsu_int8_row8_data[95]}},mxu_if.mxu_lsu_int8_row8_data[95:88]};
            tr.matrix_result_int16[8][12] = {{16{mxu_if.mxu_lsu_int16_row8_data[207]}},mxu_if.mxu_lsu_int16_row8_data[207:192]};
            tr.matrix_result_int8[8][12] = {{24{mxu_if.mxu_lsu_int8_row8_data[103]}},mxu_if.mxu_lsu_int8_row8_data[103:96]};
            tr.matrix_result_int16[8][13] = {{16{mxu_if.mxu_lsu_int16_row8_data[223]}},mxu_if.mxu_lsu_int16_row8_data[223:208]};
            tr.matrix_result_int8[8][13] = {{24{mxu_if.mxu_lsu_int8_row8_data[111]}},mxu_if.mxu_lsu_int8_row8_data[111:104]};
            tr.matrix_result_int16[8][14] = {{16{mxu_if.mxu_lsu_int16_row8_data[239]}},mxu_if.mxu_lsu_int16_row8_data[239:224]};
            tr.matrix_result_int8[8][14] = {{24{mxu_if.mxu_lsu_int8_row8_data[119]}},mxu_if.mxu_lsu_int8_row8_data[119:112]};
            tr.matrix_result_int16[8][15] = {{16{mxu_if.mxu_lsu_int16_row8_data[255]}},mxu_if.mxu_lsu_int16_row8_data[255:240]};
            tr.matrix_result_int8[8][15] = {{24{mxu_if.mxu_lsu_int8_row8_data[127]}},mxu_if.mxu_lsu_int8_row8_data[127:120]};
            tr.matrix_result_int16[9][0] = {{16{mxu_if.mxu_lsu_int16_row9_data[15]}},mxu_if.mxu_lsu_int16_row9_data[15:0]};
            tr.matrix_result_int8[9][0] = {{24{mxu_if.mxu_lsu_int8_row9_data[7]}},mxu_if.mxu_lsu_int8_row9_data[7:0]};
            tr.matrix_result_int16[9][1] = {{16{mxu_if.mxu_lsu_int16_row9_data[31]}},mxu_if.mxu_lsu_int16_row9_data[31:16]};
            tr.matrix_result_int8[9][1] = {{24{mxu_if.mxu_lsu_int8_row9_data[15]}},mxu_if.mxu_lsu_int8_row9_data[15:8]};
            tr.matrix_result_int16[9][2] = {{16{mxu_if.mxu_lsu_int16_row9_data[47]}},mxu_if.mxu_lsu_int16_row9_data[47:32]};
            tr.matrix_result_int8[9][2] = {{24{mxu_if.mxu_lsu_int8_row9_data[23]}},mxu_if.mxu_lsu_int8_row9_data[23:16]};
            tr.matrix_result_int16[9][3] = {{16{mxu_if.mxu_lsu_int16_row9_data[63]}},mxu_if.mxu_lsu_int16_row9_data[63:48]};
            tr.matrix_result_int8[9][3] = {{24{mxu_if.mxu_lsu_int8_row9_data[31]}},mxu_if.mxu_lsu_int8_row9_data[31:24]};
            tr.matrix_result_int16[9][4] = {{16{mxu_if.mxu_lsu_int16_row9_data[79]}},mxu_if.mxu_lsu_int16_row9_data[79:64]};
            tr.matrix_result_int8[9][4] = {{24{mxu_if.mxu_lsu_int8_row9_data[39]}},mxu_if.mxu_lsu_int8_row9_data[39:32]};
            tr.matrix_result_int16[9][5] = {{16{mxu_if.mxu_lsu_int16_row9_data[95]}},mxu_if.mxu_lsu_int16_row9_data[95:80]};
            tr.matrix_result_int8[9][5] = {{24{mxu_if.mxu_lsu_int8_row9_data[47]}},mxu_if.mxu_lsu_int8_row9_data[47:40]};
            tr.matrix_result_int16[9][6] = {{16{mxu_if.mxu_lsu_int16_row9_data[111]}},mxu_if.mxu_lsu_int16_row9_data[111:96]};
            tr.matrix_result_int8[9][6] = {{24{mxu_if.mxu_lsu_int8_row9_data[55]}},mxu_if.mxu_lsu_int8_row9_data[55:48]};
            tr.matrix_result_int16[9][7] = {{16{mxu_if.mxu_lsu_int16_row9_data[127]}},mxu_if.mxu_lsu_int16_row9_data[127:112]};
            tr.matrix_result_int8[9][7] = {{24{mxu_if.mxu_lsu_int8_row9_data[63]}},mxu_if.mxu_lsu_int8_row9_data[63:56]};
            tr.matrix_result_int16[9][8] = {{16{mxu_if.mxu_lsu_int16_row9_data[143]}},mxu_if.mxu_lsu_int16_row9_data[143:128]};
            tr.matrix_result_int8[9][8] = {{24{mxu_if.mxu_lsu_int8_row9_data[71]}},mxu_if.mxu_lsu_int8_row9_data[71:64]};
            tr.matrix_result_int16[9][9] = {{16{mxu_if.mxu_lsu_int16_row9_data[159]}},mxu_if.mxu_lsu_int16_row9_data[159:144]};
            tr.matrix_result_int8[9][9] = {{24{mxu_if.mxu_lsu_int8_row9_data[79]}},mxu_if.mxu_lsu_int8_row9_data[79:72]};
            tr.matrix_result_int16[9][10] = {{16{mxu_if.mxu_lsu_int16_row9_data[175]}},mxu_if.mxu_lsu_int16_row9_data[175:160]};
            tr.matrix_result_int8[9][10] = {{24{mxu_if.mxu_lsu_int8_row9_data[87]}},mxu_if.mxu_lsu_int8_row9_data[87:80]};
            tr.matrix_result_int16[9][11] = {{16{mxu_if.mxu_lsu_int16_row9_data[191]}},mxu_if.mxu_lsu_int16_row9_data[191:176]};
            tr.matrix_result_int8[9][11] = {{24{mxu_if.mxu_lsu_int8_row9_data[95]}},mxu_if.mxu_lsu_int8_row9_data[95:88]};
            tr.matrix_result_int16[9][12] = {{16{mxu_if.mxu_lsu_int16_row9_data[207]}},mxu_if.mxu_lsu_int16_row9_data[207:192]};
            tr.matrix_result_int8[9][12] = {{24{mxu_if.mxu_lsu_int8_row9_data[103]}},mxu_if.mxu_lsu_int8_row9_data[103:96]};
            tr.matrix_result_int16[9][13] = {{16{mxu_if.mxu_lsu_int16_row9_data[223]}},mxu_if.mxu_lsu_int16_row9_data[223:208]};
            tr.matrix_result_int8[9][13] = {{24{mxu_if.mxu_lsu_int8_row9_data[111]}},mxu_if.mxu_lsu_int8_row9_data[111:104]};
            tr.matrix_result_int16[9][14] = {{16{mxu_if.mxu_lsu_int16_row9_data[239]}},mxu_if.mxu_lsu_int16_row9_data[239:224]};
            tr.matrix_result_int8[9][14] = {{24{mxu_if.mxu_lsu_int8_row9_data[119]}},mxu_if.mxu_lsu_int8_row9_data[119:112]};
            tr.matrix_result_int16[9][15] = {{16{mxu_if.mxu_lsu_int16_row9_data[255]}},mxu_if.mxu_lsu_int16_row9_data[255:240]};
            tr.matrix_result_int8[9][15] = {{24{mxu_if.mxu_lsu_int8_row9_data[127]}},mxu_if.mxu_lsu_int8_row9_data[127:120]};
            tr.matrix_result_int16[10][0] = {{16{mxu_if.mxu_lsu_int16_row10_data[15]}},mxu_if.mxu_lsu_int16_row10_data[15:0]};
            tr.matrix_result_int8[10][0] = {{24{mxu_if.mxu_lsu_int8_row10_data[7]}},mxu_if.mxu_lsu_int8_row10_data[7:0]};
            tr.matrix_result_int16[10][1] = {{16{mxu_if.mxu_lsu_int16_row10_data[31]}},mxu_if.mxu_lsu_int16_row10_data[31:16]};
            tr.matrix_result_int8[10][1] = {{24{mxu_if.mxu_lsu_int8_row10_data[15]}},mxu_if.mxu_lsu_int8_row10_data[15:8]};
            tr.matrix_result_int16[10][2] = {{16{mxu_if.mxu_lsu_int16_row10_data[47]}},mxu_if.mxu_lsu_int16_row10_data[47:32]};
            tr.matrix_result_int8[10][2] = {{24{mxu_if.mxu_lsu_int8_row10_data[23]}},mxu_if.mxu_lsu_int8_row10_data[23:16]};
            tr.matrix_result_int16[10][3] = {{16{mxu_if.mxu_lsu_int16_row10_data[63]}},mxu_if.mxu_lsu_int16_row10_data[63:48]};
            tr.matrix_result_int8[10][3] = {{24{mxu_if.mxu_lsu_int8_row10_data[31]}},mxu_if.mxu_lsu_int8_row10_data[31:24]};
            tr.matrix_result_int16[10][4] = {{16{mxu_if.mxu_lsu_int16_row10_data[79]}},mxu_if.mxu_lsu_int16_row10_data[79:64]};
            tr.matrix_result_int8[10][4] = {{24{mxu_if.mxu_lsu_int8_row10_data[39]}},mxu_if.mxu_lsu_int8_row10_data[39:32]};
            tr.matrix_result_int16[10][5] = {{16{mxu_if.mxu_lsu_int16_row10_data[95]}},mxu_if.mxu_lsu_int16_row10_data[95:80]};
            tr.matrix_result_int8[10][5] = {{24{mxu_if.mxu_lsu_int8_row10_data[47]}},mxu_if.mxu_lsu_int8_row10_data[47:40]};
            tr.matrix_result_int16[10][6] = {{16{mxu_if.mxu_lsu_int16_row10_data[111]}},mxu_if.mxu_lsu_int16_row10_data[111:96]};
            tr.matrix_result_int8[10][6] = {{24{mxu_if.mxu_lsu_int8_row10_data[55]}},mxu_if.mxu_lsu_int8_row10_data[55:48]};
            tr.matrix_result_int16[10][7] = {{16{mxu_if.mxu_lsu_int16_row10_data[127]}},mxu_if.mxu_lsu_int16_row10_data[127:112]};
            tr.matrix_result_int8[10][7] = {{24{mxu_if.mxu_lsu_int8_row10_data[63]}},mxu_if.mxu_lsu_int8_row10_data[63:56]};
            tr.matrix_result_int16[10][8] = {{16{mxu_if.mxu_lsu_int16_row10_data[143]}},mxu_if.mxu_lsu_int16_row10_data[143:128]};
            tr.matrix_result_int8[10][8] = {{24{mxu_if.mxu_lsu_int8_row10_data[71]}},mxu_if.mxu_lsu_int8_row10_data[71:64]};
            tr.matrix_result_int16[10][9] = {{16{mxu_if.mxu_lsu_int16_row10_data[159]}},mxu_if.mxu_lsu_int16_row10_data[159:144]};
            tr.matrix_result_int8[10][9] = {{24{mxu_if.mxu_lsu_int8_row10_data[79]}},mxu_if.mxu_lsu_int8_row10_data[79:72]};
            tr.matrix_result_int16[10][10] = {{16{mxu_if.mxu_lsu_int16_row10_data[175]}},mxu_if.mxu_lsu_int16_row10_data[175:160]};
            tr.matrix_result_int8[10][10] = {{24{mxu_if.mxu_lsu_int8_row10_data[87]}},mxu_if.mxu_lsu_int8_row10_data[87:80]};
            tr.matrix_result_int16[10][11] = {{16{mxu_if.mxu_lsu_int16_row10_data[191]}},mxu_if.mxu_lsu_int16_row10_data[191:176]};
            tr.matrix_result_int8[10][11] = {{24{mxu_if.mxu_lsu_int8_row10_data[95]}},mxu_if.mxu_lsu_int8_row10_data[95:88]};
            tr.matrix_result_int16[10][12] = {{16{mxu_if.mxu_lsu_int16_row10_data[207]}},mxu_if.mxu_lsu_int16_row10_data[207:192]};
            tr.matrix_result_int8[10][12] = {{24{mxu_if.mxu_lsu_int8_row10_data[103]}},mxu_if.mxu_lsu_int8_row10_data[103:96]};
            tr.matrix_result_int16[10][13] = {{16{mxu_if.mxu_lsu_int16_row10_data[223]}},mxu_if.mxu_lsu_int16_row10_data[223:208]};
            tr.matrix_result_int8[10][13] = {{24{mxu_if.mxu_lsu_int8_row10_data[111]}},mxu_if.mxu_lsu_int8_row10_data[111:104]};
            tr.matrix_result_int16[10][14] = {{16{mxu_if.mxu_lsu_int16_row10_data[239]}},mxu_if.mxu_lsu_int16_row10_data[239:224]};
            tr.matrix_result_int8[10][14] = {{24{mxu_if.mxu_lsu_int8_row10_data[119]}},mxu_if.mxu_lsu_int8_row10_data[119:112]};
            tr.matrix_result_int16[10][15] = {{16{mxu_if.mxu_lsu_int16_row10_data[255]}},mxu_if.mxu_lsu_int16_row10_data[255:240]};
            tr.matrix_result_int8[10][15] = {{24{mxu_if.mxu_lsu_int8_row10_data[127]}},mxu_if.mxu_lsu_int8_row10_data[127:120]};
            tr.matrix_result_int16[11][0] = {{16{mxu_if.mxu_lsu_int16_row11_data[15]}},mxu_if.mxu_lsu_int16_row11_data[15:0]};
            tr.matrix_result_int8[11][0] = {{24{mxu_if.mxu_lsu_int8_row11_data[7]}},mxu_if.mxu_lsu_int8_row11_data[7:0]};
            tr.matrix_result_int16[11][1] = {{16{mxu_if.mxu_lsu_int16_row11_data[31]}},mxu_if.mxu_lsu_int16_row11_data[31:16]};
            tr.matrix_result_int8[11][1] = {{24{mxu_if.mxu_lsu_int8_row11_data[15]}},mxu_if.mxu_lsu_int8_row11_data[15:8]};
            tr.matrix_result_int16[11][2] = {{16{mxu_if.mxu_lsu_int16_row11_data[47]}},mxu_if.mxu_lsu_int16_row11_data[47:32]};
            tr.matrix_result_int8[11][2] = {{24{mxu_if.mxu_lsu_int8_row11_data[23]}},mxu_if.mxu_lsu_int8_row11_data[23:16]};
            tr.matrix_result_int16[11][3] = {{16{mxu_if.mxu_lsu_int16_row11_data[63]}},mxu_if.mxu_lsu_int16_row11_data[63:48]};
            tr.matrix_result_int8[11][3] = {{24{mxu_if.mxu_lsu_int8_row11_data[31]}},mxu_if.mxu_lsu_int8_row11_data[31:24]};
            tr.matrix_result_int16[11][4] = {{16{mxu_if.mxu_lsu_int16_row11_data[79]}},mxu_if.mxu_lsu_int16_row11_data[79:64]};
            tr.matrix_result_int8[11][4] = {{24{mxu_if.mxu_lsu_int8_row11_data[39]}},mxu_if.mxu_lsu_int8_row11_data[39:32]};
            tr.matrix_result_int16[11][5] = {{16{mxu_if.mxu_lsu_int16_row11_data[95]}},mxu_if.mxu_lsu_int16_row11_data[95:80]};
            tr.matrix_result_int8[11][5] = {{24{mxu_if.mxu_lsu_int8_row11_data[47]}},mxu_if.mxu_lsu_int8_row11_data[47:40]};
            tr.matrix_result_int16[11][6] = {{16{mxu_if.mxu_lsu_int16_row11_data[111]}},mxu_if.mxu_lsu_int16_row11_data[111:96]};
            tr.matrix_result_int8[11][6] = {{24{mxu_if.mxu_lsu_int8_row11_data[55]}},mxu_if.mxu_lsu_int8_row11_data[55:48]};
            tr.matrix_result_int16[11][7] = {{16{mxu_if.mxu_lsu_int16_row11_data[127]}},mxu_if.mxu_lsu_int16_row11_data[127:112]};
            tr.matrix_result_int8[11][7] = {{24{mxu_if.mxu_lsu_int8_row11_data[63]}},mxu_if.mxu_lsu_int8_row11_data[63:56]};
            tr.matrix_result_int16[11][8] = {{16{mxu_if.mxu_lsu_int16_row11_data[143]}},mxu_if.mxu_lsu_int16_row11_data[143:128]};
            tr.matrix_result_int8[11][8] = {{24{mxu_if.mxu_lsu_int8_row11_data[71]}},mxu_if.mxu_lsu_int8_row11_data[71:64]};
            tr.matrix_result_int16[11][9] = {{16{mxu_if.mxu_lsu_int16_row11_data[159]}},mxu_if.mxu_lsu_int16_row11_data[159:144]};
            tr.matrix_result_int8[11][9] = {{24{mxu_if.mxu_lsu_int8_row11_data[79]}},mxu_if.mxu_lsu_int8_row11_data[79:72]};
            tr.matrix_result_int16[11][10] = {{16{mxu_if.mxu_lsu_int16_row11_data[175]}},mxu_if.mxu_lsu_int16_row11_data[175:160]};
            tr.matrix_result_int8[11][10] = {{24{mxu_if.mxu_lsu_int8_row11_data[87]}},mxu_if.mxu_lsu_int8_row11_data[87:80]};
            tr.matrix_result_int16[11][11] = {{16{mxu_if.mxu_lsu_int16_row11_data[191]}},mxu_if.mxu_lsu_int16_row11_data[191:176]};
            tr.matrix_result_int8[11][11] = {{24{mxu_if.mxu_lsu_int8_row11_data[95]}},mxu_if.mxu_lsu_int8_row11_data[95:88]};
            tr.matrix_result_int16[11][12] = {{16{mxu_if.mxu_lsu_int16_row11_data[207]}},mxu_if.mxu_lsu_int16_row11_data[207:192]};
            tr.matrix_result_int8[11][12] = {{24{mxu_if.mxu_lsu_int8_row11_data[103]}},mxu_if.mxu_lsu_int8_row11_data[103:96]};
            tr.matrix_result_int16[11][13] = {{16{mxu_if.mxu_lsu_int16_row11_data[223]}},mxu_if.mxu_lsu_int16_row11_data[223:208]};
            tr.matrix_result_int8[11][13] = {{24{mxu_if.mxu_lsu_int8_row11_data[111]}},mxu_if.mxu_lsu_int8_row11_data[111:104]};
            tr.matrix_result_int16[11][14] = {{16{mxu_if.mxu_lsu_int16_row11_data[239]}},mxu_if.mxu_lsu_int16_row11_data[239:224]};
            tr.matrix_result_int8[11][14] = {{24{mxu_if.mxu_lsu_int8_row11_data[119]}},mxu_if.mxu_lsu_int8_row11_data[119:112]};
            tr.matrix_result_int16[11][15] = {{16{mxu_if.mxu_lsu_int16_row11_data[255]}},mxu_if.mxu_lsu_int16_row11_data[255:240]};
            tr.matrix_result_int8[11][15] = {{24{mxu_if.mxu_lsu_int8_row11_data[127]}},mxu_if.mxu_lsu_int8_row11_data[127:120]};
            tr.matrix_result_int16[12][0] = {{16{mxu_if.mxu_lsu_int16_row12_data[15]}},mxu_if.mxu_lsu_int16_row12_data[15:0]};
            tr.matrix_result_int8[12][0] = {{24{mxu_if.mxu_lsu_int8_row12_data[7]}},mxu_if.mxu_lsu_int8_row12_data[7:0]};
            tr.matrix_result_int16[12][1] = {{16{mxu_if.mxu_lsu_int16_row12_data[31]}},mxu_if.mxu_lsu_int16_row12_data[31:16]};
            tr.matrix_result_int8[12][1] = {{24{mxu_if.mxu_lsu_int8_row12_data[15]}},mxu_if.mxu_lsu_int8_row12_data[15:8]};
            tr.matrix_result_int16[12][2] = {{16{mxu_if.mxu_lsu_int16_row12_data[47]}},mxu_if.mxu_lsu_int16_row12_data[47:32]};
            tr.matrix_result_int8[12][2] = {{24{mxu_if.mxu_lsu_int8_row12_data[23]}},mxu_if.mxu_lsu_int8_row12_data[23:16]};
            tr.matrix_result_int16[12][3] = {{16{mxu_if.mxu_lsu_int16_row12_data[63]}},mxu_if.mxu_lsu_int16_row12_data[63:48]};
            tr.matrix_result_int8[12][3] = {{24{mxu_if.mxu_lsu_int8_row12_data[31]}},mxu_if.mxu_lsu_int8_row12_data[31:24]};
            tr.matrix_result_int16[12][4] = {{16{mxu_if.mxu_lsu_int16_row12_data[79]}},mxu_if.mxu_lsu_int16_row12_data[79:64]};
            tr.matrix_result_int8[12][4] = {{24{mxu_if.mxu_lsu_int8_row12_data[39]}},mxu_if.mxu_lsu_int8_row12_data[39:32]};
            tr.matrix_result_int16[12][5] = {{16{mxu_if.mxu_lsu_int16_row12_data[95]}},mxu_if.mxu_lsu_int16_row12_data[95:80]};
            tr.matrix_result_int8[12][5] = {{24{mxu_if.mxu_lsu_int8_row12_data[47]}},mxu_if.mxu_lsu_int8_row12_data[47:40]};
            tr.matrix_result_int16[12][6] = {{16{mxu_if.mxu_lsu_int16_row12_data[111]}},mxu_if.mxu_lsu_int16_row12_data[111:96]};
            tr.matrix_result_int8[12][6] = {{24{mxu_if.mxu_lsu_int8_row12_data[55]}},mxu_if.mxu_lsu_int8_row12_data[55:48]};
            tr.matrix_result_int16[12][7] = {{16{mxu_if.mxu_lsu_int16_row12_data[127]}},mxu_if.mxu_lsu_int16_row12_data[127:112]};
            tr.matrix_result_int8[12][7] = {{24{mxu_if.mxu_lsu_int8_row12_data[63]}},mxu_if.mxu_lsu_int8_row12_data[63:56]};
            tr.matrix_result_int16[12][8] = {{16{mxu_if.mxu_lsu_int16_row12_data[143]}},mxu_if.mxu_lsu_int16_row12_data[143:128]};
            tr.matrix_result_int8[12][8] = {{24{mxu_if.mxu_lsu_int8_row12_data[71]}},mxu_if.mxu_lsu_int8_row12_data[71:64]};
            tr.matrix_result_int16[12][9] = {{16{mxu_if.mxu_lsu_int16_row12_data[159]}},mxu_if.mxu_lsu_int16_row12_data[159:144]};
            tr.matrix_result_int8[12][9] = {{24{mxu_if.mxu_lsu_int8_row12_data[79]}},mxu_if.mxu_lsu_int8_row12_data[79:72]};
            tr.matrix_result_int16[12][10] = {{16{mxu_if.mxu_lsu_int16_row12_data[175]}},mxu_if.mxu_lsu_int16_row12_data[175:160]};
            tr.matrix_result_int8[12][10] = {{24{mxu_if.mxu_lsu_int8_row12_data[87]}},mxu_if.mxu_lsu_int8_row12_data[87:80]};
            tr.matrix_result_int16[12][11] = {{16{mxu_if.mxu_lsu_int16_row12_data[191]}},mxu_if.mxu_lsu_int16_row12_data[191:176]};
            tr.matrix_result_int8[12][11] = {{24{mxu_if.mxu_lsu_int8_row12_data[95]}},mxu_if.mxu_lsu_int8_row12_data[95:88]};
            tr.matrix_result_int16[12][12] = {{16{mxu_if.mxu_lsu_int16_row12_data[207]}},mxu_if.mxu_lsu_int16_row12_data[207:192]};
            tr.matrix_result_int8[12][12] = {{24{mxu_if.mxu_lsu_int8_row12_data[103]}},mxu_if.mxu_lsu_int8_row12_data[103:96]};
            tr.matrix_result_int16[12][13] = {{16{mxu_if.mxu_lsu_int16_row12_data[223]}},mxu_if.mxu_lsu_int16_row12_data[223:208]};
            tr.matrix_result_int8[12][13] = {{24{mxu_if.mxu_lsu_int8_row12_data[111]}},mxu_if.mxu_lsu_int8_row12_data[111:104]};
            tr.matrix_result_int16[12][14] = {{16{mxu_if.mxu_lsu_int16_row12_data[239]}},mxu_if.mxu_lsu_int16_row12_data[239:224]};
            tr.matrix_result_int8[12][14] = {{24{mxu_if.mxu_lsu_int8_row12_data[119]}},mxu_if.mxu_lsu_int8_row12_data[119:112]};
            tr.matrix_result_int16[12][15] = {{16{mxu_if.mxu_lsu_int16_row12_data[255]}},mxu_if.mxu_lsu_int16_row12_data[255:240]};
            tr.matrix_result_int8[12][15] = {{24{mxu_if.mxu_lsu_int8_row12_data[127]}},mxu_if.mxu_lsu_int8_row12_data[127:120]};
            tr.matrix_result_int16[13][0] = {{16{mxu_if.mxu_lsu_int16_row13_data[15]}},mxu_if.mxu_lsu_int16_row13_data[15:0]};
            tr.matrix_result_int8[13][0] = {{24{mxu_if.mxu_lsu_int8_row13_data[7]}},mxu_if.mxu_lsu_int8_row13_data[7:0]};
            tr.matrix_result_int16[13][1] = {{16{mxu_if.mxu_lsu_int16_row13_data[31]}},mxu_if.mxu_lsu_int16_row13_data[31:16]};
            tr.matrix_result_int8[13][1] = {{24{mxu_if.mxu_lsu_int8_row13_data[15]}},mxu_if.mxu_lsu_int8_row13_data[15:8]};
            tr.matrix_result_int16[13][2] = {{16{mxu_if.mxu_lsu_int16_row13_data[47]}},mxu_if.mxu_lsu_int16_row13_data[47:32]};
            tr.matrix_result_int8[13][2] = {{24{mxu_if.mxu_lsu_int8_row13_data[23]}},mxu_if.mxu_lsu_int8_row13_data[23:16]};
            tr.matrix_result_int16[13][3] = {{16{mxu_if.mxu_lsu_int16_row13_data[63]}},mxu_if.mxu_lsu_int16_row13_data[63:48]};
            tr.matrix_result_int8[13][3] = {{24{mxu_if.mxu_lsu_int8_row13_data[31]}},mxu_if.mxu_lsu_int8_row13_data[31:24]};
            tr.matrix_result_int16[13][4] = {{16{mxu_if.mxu_lsu_int16_row13_data[79]}},mxu_if.mxu_lsu_int16_row13_data[79:64]};
            tr.matrix_result_int8[13][4] = {{24{mxu_if.mxu_lsu_int8_row13_data[39]}},mxu_if.mxu_lsu_int8_row13_data[39:32]};
            tr.matrix_result_int16[13][5] = {{16{mxu_if.mxu_lsu_int16_row13_data[95]}},mxu_if.mxu_lsu_int16_row13_data[95:80]};
            tr.matrix_result_int8[13][5] = {{24{mxu_if.mxu_lsu_int8_row13_data[47]}},mxu_if.mxu_lsu_int8_row13_data[47:40]};
            tr.matrix_result_int16[13][6] = {{16{mxu_if.mxu_lsu_int16_row13_data[111]}},mxu_if.mxu_lsu_int16_row13_data[111:96]};
            tr.matrix_result_int8[13][6] = {{24{mxu_if.mxu_lsu_int8_row13_data[55]}},mxu_if.mxu_lsu_int8_row13_data[55:48]};
            tr.matrix_result_int16[13][7] = {{16{mxu_if.mxu_lsu_int16_row13_data[127]}},mxu_if.mxu_lsu_int16_row13_data[127:112]};
            tr.matrix_result_int8[13][7] = {{24{mxu_if.mxu_lsu_int8_row13_data[63]}},mxu_if.mxu_lsu_int8_row13_data[63:56]};
            tr.matrix_result_int16[13][8] = {{16{mxu_if.mxu_lsu_int16_row13_data[143]}},mxu_if.mxu_lsu_int16_row13_data[143:128]};
            tr.matrix_result_int8[13][8] = {{24{mxu_if.mxu_lsu_int8_row13_data[71]}},mxu_if.mxu_lsu_int8_row13_data[71:64]};
            tr.matrix_result_int16[13][9] = {{16{mxu_if.mxu_lsu_int16_row13_data[159]}},mxu_if.mxu_lsu_int16_row13_data[159:144]};
            tr.matrix_result_int8[13][9] = {{24{mxu_if.mxu_lsu_int8_row13_data[79]}},mxu_if.mxu_lsu_int8_row13_data[79:72]};
            tr.matrix_result_int16[13][10] = {{16{mxu_if.mxu_lsu_int16_row13_data[175]}},mxu_if.mxu_lsu_int16_row13_data[175:160]};
            tr.matrix_result_int8[13][10] = {{24{mxu_if.mxu_lsu_int8_row13_data[87]}},mxu_if.mxu_lsu_int8_row13_data[87:80]};
            tr.matrix_result_int16[13][11] = {{16{mxu_if.mxu_lsu_int16_row13_data[191]}},mxu_if.mxu_lsu_int16_row13_data[191:176]};
            tr.matrix_result_int8[13][11] = {{24{mxu_if.mxu_lsu_int8_row13_data[95]}},mxu_if.mxu_lsu_int8_row13_data[95:88]};
            tr.matrix_result_int16[13][12] = {{16{mxu_if.mxu_lsu_int16_row13_data[207]}},mxu_if.mxu_lsu_int16_row13_data[207:192]};
            tr.matrix_result_int8[13][12] = {{24{mxu_if.mxu_lsu_int8_row13_data[103]}},mxu_if.mxu_lsu_int8_row13_data[103:96]};
            tr.matrix_result_int16[13][13] = {{16{mxu_if.mxu_lsu_int16_row13_data[223]}},mxu_if.mxu_lsu_int16_row13_data[223:208]};
            tr.matrix_result_int8[13][13] = {{24{mxu_if.mxu_lsu_int8_row13_data[111]}},mxu_if.mxu_lsu_int8_row13_data[111:104]};
            tr.matrix_result_int16[13][14] = {{16{mxu_if.mxu_lsu_int16_row13_data[239]}},mxu_if.mxu_lsu_int16_row13_data[239:224]};
            tr.matrix_result_int8[13][14] = {{24{mxu_if.mxu_lsu_int8_row13_data[119]}},mxu_if.mxu_lsu_int8_row13_data[119:112]};
            tr.matrix_result_int16[13][15] = {{16{mxu_if.mxu_lsu_int16_row13_data[255]}},mxu_if.mxu_lsu_int16_row13_data[255:240]};
            tr.matrix_result_int8[13][15] = {{24{mxu_if.mxu_lsu_int8_row13_data[127]}},mxu_if.mxu_lsu_int8_row13_data[127:120]};
            tr.matrix_result_int16[14][0] = {{16{mxu_if.mxu_lsu_int16_row14_data[15]}},mxu_if.mxu_lsu_int16_row14_data[15:0]};
            tr.matrix_result_int8[14][0] = {{24{mxu_if.mxu_lsu_int8_row14_data[7]}},mxu_if.mxu_lsu_int8_row14_data[7:0]};
            tr.matrix_result_int16[14][1] = {{16{mxu_if.mxu_lsu_int16_row14_data[31]}},mxu_if.mxu_lsu_int16_row14_data[31:16]};
            tr.matrix_result_int8[14][1] = {{24{mxu_if.mxu_lsu_int8_row14_data[15]}},mxu_if.mxu_lsu_int8_row14_data[15:8]};
            tr.matrix_result_int16[14][2] = {{16{mxu_if.mxu_lsu_int16_row14_data[47]}},mxu_if.mxu_lsu_int16_row14_data[47:32]};
            tr.matrix_result_int8[14][2] = {{24{mxu_if.mxu_lsu_int8_row14_data[23]}},mxu_if.mxu_lsu_int8_row14_data[23:16]};
            tr.matrix_result_int16[14][3] = {{16{mxu_if.mxu_lsu_int16_row14_data[63]}},mxu_if.mxu_lsu_int16_row14_data[63:48]};
            tr.matrix_result_int8[14][3] = {{24{mxu_if.mxu_lsu_int8_row14_data[31]}},mxu_if.mxu_lsu_int8_row14_data[31:24]};
            tr.matrix_result_int16[14][4] = {{16{mxu_if.mxu_lsu_int16_row14_data[79]}},mxu_if.mxu_lsu_int16_row14_data[79:64]};
            tr.matrix_result_int8[14][4] = {{24{mxu_if.mxu_lsu_int8_row14_data[39]}},mxu_if.mxu_lsu_int8_row14_data[39:32]};
            tr.matrix_result_int16[14][5] = {{16{mxu_if.mxu_lsu_int16_row14_data[95]}},mxu_if.mxu_lsu_int16_row14_data[95:80]};
            tr.matrix_result_int8[14][5] = {{24{mxu_if.mxu_lsu_int8_row14_data[47]}},mxu_if.mxu_lsu_int8_row14_data[47:40]};
            tr.matrix_result_int16[14][6] = {{16{mxu_if.mxu_lsu_int16_row14_data[111]}},mxu_if.mxu_lsu_int16_row14_data[111:96]};
            tr.matrix_result_int8[14][6] = {{24{mxu_if.mxu_lsu_int8_row14_data[55]}},mxu_if.mxu_lsu_int8_row14_data[55:48]};
            tr.matrix_result_int16[14][7] = {{16{mxu_if.mxu_lsu_int16_row14_data[127]}},mxu_if.mxu_lsu_int16_row14_data[127:112]};
            tr.matrix_result_int8[14][7] = {{24{mxu_if.mxu_lsu_int8_row14_data[63]}},mxu_if.mxu_lsu_int8_row14_data[63:56]};
            tr.matrix_result_int16[14][8] = {{16{mxu_if.mxu_lsu_int16_row14_data[143]}},mxu_if.mxu_lsu_int16_row14_data[143:128]};
            tr.matrix_result_int8[14][8] = {{24{mxu_if.mxu_lsu_int8_row14_data[71]}},mxu_if.mxu_lsu_int8_row14_data[71:64]};
            tr.matrix_result_int16[14][9] = {{16{mxu_if.mxu_lsu_int16_row14_data[159]}},mxu_if.mxu_lsu_int16_row14_data[159:144]};
            tr.matrix_result_int8[14][9] = {{24{mxu_if.mxu_lsu_int8_row14_data[79]}},mxu_if.mxu_lsu_int8_row14_data[79:72]};
            tr.matrix_result_int16[14][10] = {{16{mxu_if.mxu_lsu_int16_row14_data[175]}},mxu_if.mxu_lsu_int16_row14_data[175:160]};
            tr.matrix_result_int8[14][10] = {{24{mxu_if.mxu_lsu_int8_row14_data[87]}},mxu_if.mxu_lsu_int8_row14_data[87:80]};
            tr.matrix_result_int16[14][11] = {{16{mxu_if.mxu_lsu_int16_row14_data[191]}},mxu_if.mxu_lsu_int16_row14_data[191:176]};
            tr.matrix_result_int8[14][11] = {{24{mxu_if.mxu_lsu_int8_row14_data[95]}},mxu_if.mxu_lsu_int8_row14_data[95:88]};
            tr.matrix_result_int16[14][12] = {{16{mxu_if.mxu_lsu_int16_row14_data[207]}},mxu_if.mxu_lsu_int16_row14_data[207:192]};
            tr.matrix_result_int8[14][12] = {{24{mxu_if.mxu_lsu_int8_row14_data[103]}},mxu_if.mxu_lsu_int8_row14_data[103:96]};
            tr.matrix_result_int16[14][13] = {{16{mxu_if.mxu_lsu_int16_row14_data[223]}},mxu_if.mxu_lsu_int16_row14_data[223:208]};
            tr.matrix_result_int8[14][13] = {{24{mxu_if.mxu_lsu_int8_row14_data[111]}},mxu_if.mxu_lsu_int8_row14_data[111:104]};
            tr.matrix_result_int16[14][14] = {{16{mxu_if.mxu_lsu_int16_row14_data[239]}},mxu_if.mxu_lsu_int16_row14_data[239:224]};
            tr.matrix_result_int8[14][14] = {{24{mxu_if.mxu_lsu_int8_row14_data[119]}},mxu_if.mxu_lsu_int8_row14_data[119:112]};
            tr.matrix_result_int16[14][15] = {{16{mxu_if.mxu_lsu_int16_row14_data[255]}},mxu_if.mxu_lsu_int16_row14_data[255:240]};
            tr.matrix_result_int8[14][15] = {{24{mxu_if.mxu_lsu_int8_row14_data[127]}},mxu_if.mxu_lsu_int8_row14_data[127:120]};
            tr.matrix_result_int16[15][0] = {{16{mxu_if.mxu_lsu_int16_row15_data[15]}},mxu_if.mxu_lsu_int16_row15_data[15:0]};
            tr.matrix_result_int8[15][0] = {{24{mxu_if.mxu_lsu_int8_row15_data[7]}},mxu_if.mxu_lsu_int8_row15_data[7:0]};
            tr.matrix_result_int16[15][1] = {{16{mxu_if.mxu_lsu_int16_row15_data[31]}},mxu_if.mxu_lsu_int16_row15_data[31:16]};
            tr.matrix_result_int8[15][1] = {{24{mxu_if.mxu_lsu_int8_row15_data[15]}},mxu_if.mxu_lsu_int8_row15_data[15:8]};
            tr.matrix_result_int16[15][2] = {{16{mxu_if.mxu_lsu_int16_row15_data[47]}},mxu_if.mxu_lsu_int16_row15_data[47:32]};
            tr.matrix_result_int8[15][2] = {{24{mxu_if.mxu_lsu_int8_row15_data[23]}},mxu_if.mxu_lsu_int8_row15_data[23:16]};
            tr.matrix_result_int16[15][3] = {{16{mxu_if.mxu_lsu_int16_row15_data[63]}},mxu_if.mxu_lsu_int16_row15_data[63:48]};
            tr.matrix_result_int8[15][3] = {{24{mxu_if.mxu_lsu_int8_row15_data[31]}},mxu_if.mxu_lsu_int8_row15_data[31:24]};
            tr.matrix_result_int16[15][4] = {{16{mxu_if.mxu_lsu_int16_row15_data[79]}},mxu_if.mxu_lsu_int16_row15_data[79:64]};
            tr.matrix_result_int8[15][4] = {{24{mxu_if.mxu_lsu_int8_row15_data[39]}},mxu_if.mxu_lsu_int8_row15_data[39:32]};
            tr.matrix_result_int16[15][5] = {{16{mxu_if.mxu_lsu_int16_row15_data[95]}},mxu_if.mxu_lsu_int16_row15_data[95:80]};
            tr.matrix_result_int8[15][5] = {{24{mxu_if.mxu_lsu_int8_row15_data[47]}},mxu_if.mxu_lsu_int8_row15_data[47:40]};
            tr.matrix_result_int16[15][6] = {{16{mxu_if.mxu_lsu_int16_row15_data[111]}},mxu_if.mxu_lsu_int16_row15_data[111:96]};
            tr.matrix_result_int8[15][6] = {{24{mxu_if.mxu_lsu_int8_row15_data[55]}},mxu_if.mxu_lsu_int8_row15_data[55:48]};
            tr.matrix_result_int16[15][7] = {{16{mxu_if.mxu_lsu_int16_row15_data[127]}},mxu_if.mxu_lsu_int16_row15_data[127:112]};
            tr.matrix_result_int8[15][7] = {{24{mxu_if.mxu_lsu_int8_row15_data[63]}},mxu_if.mxu_lsu_int8_row15_data[63:56]};
            tr.matrix_result_int16[15][8] = {{16{mxu_if.mxu_lsu_int16_row15_data[143]}},mxu_if.mxu_lsu_int16_row15_data[143:128]};
            tr.matrix_result_int8[15][8] = {{24{mxu_if.mxu_lsu_int8_row15_data[71]}},mxu_if.mxu_lsu_int8_row15_data[71:64]};
            tr.matrix_result_int16[15][9] = {{16{mxu_if.mxu_lsu_int16_row15_data[159]}},mxu_if.mxu_lsu_int16_row15_data[159:144]};
            tr.matrix_result_int8[15][9] = {{24{mxu_if.mxu_lsu_int8_row15_data[79]}},mxu_if.mxu_lsu_int8_row15_data[79:72]};
            tr.matrix_result_int16[15][10] = {{16{mxu_if.mxu_lsu_int16_row15_data[175]}},mxu_if.mxu_lsu_int16_row15_data[175:160]};
            tr.matrix_result_int8[15][10] = {{24{mxu_if.mxu_lsu_int8_row15_data[87]}},mxu_if.mxu_lsu_int8_row15_data[87:80]};
            tr.matrix_result_int16[15][11] = {{16{mxu_if.mxu_lsu_int16_row15_data[191]}},mxu_if.mxu_lsu_int16_row15_data[191:176]};
            tr.matrix_result_int8[15][11] = {{24{mxu_if.mxu_lsu_int8_row15_data[95]}},mxu_if.mxu_lsu_int8_row15_data[95:88]};
            tr.matrix_result_int16[15][12] = {{16{mxu_if.mxu_lsu_int16_row15_data[207]}},mxu_if.mxu_lsu_int16_row15_data[207:192]};
            tr.matrix_result_int8[15][12] = {{24{mxu_if.mxu_lsu_int8_row15_data[103]}},mxu_if.mxu_lsu_int8_row15_data[103:96]};
            tr.matrix_result_int16[15][13] = {{16{mxu_if.mxu_lsu_int16_row15_data[223]}},mxu_if.mxu_lsu_int16_row15_data[223:208]};
            tr.matrix_result_int8[15][13] = {{24{mxu_if.mxu_lsu_int8_row15_data[111]}},mxu_if.mxu_lsu_int8_row15_data[111:104]};
            tr.matrix_result_int16[15][14] = {{16{mxu_if.mxu_lsu_int16_row15_data[239]}},mxu_if.mxu_lsu_int16_row15_data[239:224]};
            tr.matrix_result_int8[15][14] = {{24{mxu_if.mxu_lsu_int8_row15_data[119]}},mxu_if.mxu_lsu_int8_row15_data[119:112]};
            tr.matrix_result_int16[15][15] = {{16{mxu_if.mxu_lsu_int16_row15_data[255]}},mxu_if.mxu_lsu_int16_row15_data[255:240]};
            tr.matrix_result_int8[15][15] = {{24{mxu_if.mxu_lsu_int8_row15_data[127]}},mxu_if.mxu_lsu_int8_row15_data[127:120]};
            break;
        end
    end

endtask

function void mxu_output_monitor::final_phase(uvm_phase phase);
    super.final_phase(phase);
    `uvm_info("mxu_omon", $sformatf("enter fianl phase, mxu_omon send cnt is %d", send_cnt), UVM_LOW);
endfunction
