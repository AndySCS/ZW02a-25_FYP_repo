class mxu_output_monitor extends uvm_monitor;

    virtual mxu_intf mxu_if;
    uvm_analysis_port #(mxu_tr) ap;

    `uvm_component_utils(mxu_output_monitor)
    function new(string name = "mxu_output_monitor", uvm_component parent = null);
       super.new(name, parent);
    endfunction //new()
    
    extern virtual task build_phase(uvm_phase phase);
    extern virtual task main_phase(uvm_phase phase);
    
    extern virtual task collect_matrix_out(mxu_tr tr);

endclass //mxu_output_monitor extends superClass

task mxu_output_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual mxu_intf)::get(this, "", "mxu_if", mxu_if))begin
        `uvm_fatal("mxu_output_monitor", "mxu output_monitor fail to get mxu if")
    end
    ap = new("ap", this);
endtask

task mxu_output_monitor::main_phase(uvm_phase phase);
    mxu_tr tr;

    tr = new("tr");

    while (1) begin 
        this.collect_matrix(tr);
        ap.write(tr);
    end

endtask

task mxu_output_monitor::collect_matrix_out(mxu_tr tr);

    while(1)begin
        @(posedge mxu_if.clk);
        if(mxu_if.lsu_mxu_vld) break;
    end

    tr.clear_result();
    @(posedge mxu_if.clk);
    wait(mxu_if.mxu_lsu_data_rdy) 
    tr.matrix_result[0].q[0] = mxu_if.mxu_lsu_int16_row0_data[7:0];
    tr.matrix_result[0].q[1] = mxu_if.mxu_lsu_int16_row0_data[15:8];
    tr.matrix_result[0].q[2] = mxu_if.mxu_lsu_int16_row0_data[23:16];
    tr.matrix_result[0].q[3] = mxu_if.mxu_lsu_int16_row0_data[31:24];
    tr.matrix_result[0].q[4] = mxu_if.mxu_lsu_int16_row0_data[39:32];
    tr.matrix_result[0].q[5] = mxu_if.mxu_lsu_int16_row0_data[47:40];
    tr.matrix_result[0].q[6] = mxu_if.mxu_lsu_int16_row0_data[55:48];
    tr.matrix_result[0].q[7] = mxu_if.mxu_lsu_int16_row0_data[63:56];
    tr.matrix_result[0].q[8] = mxu_if.mxu_lsu_int16_row0_data[71:64];
    tr.matrix_result[0].q[9] = mxu_if.mxu_lsu_int16_row0_data[79:72];
    tr.matrix_result[0].q[10] = mxu_if.mxu_lsu_int16_row0_data[87:80];
    tr.matrix_result[0].q[11] = mxu_if.mxu_lsu_int16_row0_data[95:88];
    tr.matrix_result[0].q[12] = mxu_if.mxu_lsu_int16_row0_data[103:96];
    tr.matrix_result[0].q[13] = mxu_if.mxu_lsu_int16_row0_data[111:104];
    tr.matrix_result[0].q[14] = mxu_if.mxu_lsu_int16_row0_data[119:112];
    tr.matrix_result[0].q[15] = mxu_if.mxu_lsu_int16_row0_data[127:120];
    tr.matrix_result[1].q[0] = mxu_if.mxu_lsu_int16_row1_data[7:0];
    tr.matrix_result[1].q[1] = mxu_if.mxu_lsu_int16_row1_data[15:8];
    tr.matrix_result[1].q[2] = mxu_if.mxu_lsu_int16_row1_data[23:16];
    tr.matrix_result[1].q[3] = mxu_if.mxu_lsu_int16_row1_data[31:24];
    tr.matrix_result[1].q[4] = mxu_if.mxu_lsu_int16_row1_data[39:32];
    tr.matrix_result[1].q[5] = mxu_if.mxu_lsu_int16_row1_data[47:40];
    tr.matrix_result[1].q[6] = mxu_if.mxu_lsu_int16_row1_data[55:48];
    tr.matrix_result[1].q[7] = mxu_if.mxu_lsu_int16_row1_data[63:56];
    tr.matrix_result[1].q[8] = mxu_if.mxu_lsu_int16_row1_data[71:64];
    tr.matrix_result[1].q[9] = mxu_if.mxu_lsu_int16_row1_data[79:72];
    tr.matrix_result[1].q[10] = mxu_if.mxu_lsu_int16_row1_data[87:80];
    tr.matrix_result[1].q[11] = mxu_if.mxu_lsu_int16_row1_data[95:88];
    tr.matrix_result[1].q[12] = mxu_if.mxu_lsu_int16_row1_data[103:96];
    tr.matrix_result[1].q[13] = mxu_if.mxu_lsu_int16_row1_data[111:104];
    tr.matrix_result[1].q[14] = mxu_if.mxu_lsu_int16_row1_data[119:112];
    tr.matrix_result[1].q[15] = mxu_if.mxu_lsu_int16_row1_data[127:120];
    tr.matrix_result[2].q[0] = mxu_if.mxu_lsu_int16_row2_data[7:0];
    tr.matrix_result[2].q[1] = mxu_if.mxu_lsu_int16_row2_data[15:8];
    tr.matrix_result[2].q[2] = mxu_if.mxu_lsu_int16_row2_data[23:16];
    tr.matrix_result[2].q[3] = mxu_if.mxu_lsu_int16_row2_data[31:24];
    tr.matrix_result[2].q[4] = mxu_if.mxu_lsu_int16_row2_data[39:32];
    tr.matrix_result[2].q[5] = mxu_if.mxu_lsu_int16_row2_data[47:40];
    tr.matrix_result[2].q[6] = mxu_if.mxu_lsu_int16_row2_data[55:48];
    tr.matrix_result[2].q[7] = mxu_if.mxu_lsu_int16_row2_data[63:56];
    tr.matrix_result[2].q[8] = mxu_if.mxu_lsu_int16_row2_data[71:64];
    tr.matrix_result[2].q[9] = mxu_if.mxu_lsu_int16_row2_data[79:72];
    tr.matrix_result[2].q[10] = mxu_if.mxu_lsu_int16_row2_data[87:80];
    tr.matrix_result[2].q[11] = mxu_if.mxu_lsu_int16_row2_data[95:88];
    tr.matrix_result[2].q[12] = mxu_if.mxu_lsu_int16_row2_data[103:96];
    tr.matrix_result[2].q[13] = mxu_if.mxu_lsu_int16_row2_data[111:104];
    tr.matrix_result[2].q[14] = mxu_if.mxu_lsu_int16_row2_data[119:112];
    tr.matrix_result[2].q[15] = mxu_if.mxu_lsu_int16_row2_data[127:120];
    tr.matrix_result[3].q[0] = mxu_if.mxu_lsu_int16_row3_data[7:0];
    tr.matrix_result[3].q[1] = mxu_if.mxu_lsu_int16_row3_data[15:8];
    tr.matrix_result[3].q[2] = mxu_if.mxu_lsu_int16_row3_data[23:16];
    tr.matrix_result[3].q[3] = mxu_if.mxu_lsu_int16_row3_data[31:24];
    tr.matrix_result[3].q[4] = mxu_if.mxu_lsu_int16_row3_data[39:32];
    tr.matrix_result[3].q[5] = mxu_if.mxu_lsu_int16_row3_data[47:40];
    tr.matrix_result[3].q[6] = mxu_if.mxu_lsu_int16_row3_data[55:48];
    tr.matrix_result[3].q[7] = mxu_if.mxu_lsu_int16_row3_data[63:56];
    tr.matrix_result[3].q[8] = mxu_if.mxu_lsu_int16_row3_data[71:64];
    tr.matrix_result[3].q[9] = mxu_if.mxu_lsu_int16_row3_data[79:72];
    tr.matrix_result[3].q[10] = mxu_if.mxu_lsu_int16_row3_data[87:80];
    tr.matrix_result[3].q[11] = mxu_if.mxu_lsu_int16_row3_data[95:88];
    tr.matrix_result[3].q[12] = mxu_if.mxu_lsu_int16_row3_data[103:96];
    tr.matrix_result[3].q[13] = mxu_if.mxu_lsu_int16_row3_data[111:104];
    tr.matrix_result[3].q[14] = mxu_if.mxu_lsu_int16_row3_data[119:112];
    tr.matrix_result[3].q[15] = mxu_if.mxu_lsu_int16_row3_data[127:120];
    tr.matrix_result[4].q[0] = mxu_if.mxu_lsu_int16_row4_data[7:0];
    tr.matrix_result[4].q[1] = mxu_if.mxu_lsu_int16_row4_data[15:8];
    tr.matrix_result[4].q[2] = mxu_if.mxu_lsu_int16_row4_data[23:16];
    tr.matrix_result[4].q[3] = mxu_if.mxu_lsu_int16_row4_data[31:24];
    tr.matrix_result[4].q[4] = mxu_if.mxu_lsu_int16_row4_data[39:32];
    tr.matrix_result[4].q[5] = mxu_if.mxu_lsu_int16_row4_data[47:40];
    tr.matrix_result[4].q[6] = mxu_if.mxu_lsu_int16_row4_data[55:48];
    tr.matrix_result[4].q[7] = mxu_if.mxu_lsu_int16_row4_data[63:56];
    tr.matrix_result[4].q[8] = mxu_if.mxu_lsu_int16_row4_data[71:64];
    tr.matrix_result[4].q[9] = mxu_if.mxu_lsu_int16_row4_data[79:72];
    tr.matrix_result[4].q[10] = mxu_if.mxu_lsu_int16_row4_data[87:80];
    tr.matrix_result[4].q[11] = mxu_if.mxu_lsu_int16_row4_data[95:88];
    tr.matrix_result[4].q[12] = mxu_if.mxu_lsu_int16_row4_data[103:96];
    tr.matrix_result[4].q[13] = mxu_if.mxu_lsu_int16_row4_data[111:104];
    tr.matrix_result[4].q[14] = mxu_if.mxu_lsu_int16_row4_data[119:112];
    tr.matrix_result[4].q[15] = mxu_if.mxu_lsu_int16_row4_data[127:120];
    tr.matrix_result[5].q[0] = mxu_if.mxu_lsu_int16_row5_data[7:0];
    tr.matrix_result[5].q[1] = mxu_if.mxu_lsu_int16_row5_data[15:8];
    tr.matrix_result[5].q[2] = mxu_if.mxu_lsu_int16_row5_data[23:16];
    tr.matrix_result[5].q[3] = mxu_if.mxu_lsu_int16_row5_data[31:24];
    tr.matrix_result[5].q[4] = mxu_if.mxu_lsu_int16_row5_data[39:32];
    tr.matrix_result[5].q[5] = mxu_if.mxu_lsu_int16_row5_data[47:40];
    tr.matrix_result[5].q[6] = mxu_if.mxu_lsu_int16_row5_data[55:48];
    tr.matrix_result[5].q[7] = mxu_if.mxu_lsu_int16_row5_data[63:56];
    tr.matrix_result[5].q[8] = mxu_if.mxu_lsu_int16_row5_data[71:64];
    tr.matrix_result[5].q[9] = mxu_if.mxu_lsu_int16_row5_data[79:72];
    tr.matrix_result[5].q[10] = mxu_if.mxu_lsu_int16_row5_data[87:80];
    tr.matrix_result[5].q[11] = mxu_if.mxu_lsu_int16_row5_data[95:88];
    tr.matrix_result[5].q[12] = mxu_if.mxu_lsu_int16_row5_data[103:96];
    tr.matrix_result[5].q[13] = mxu_if.mxu_lsu_int16_row5_data[111:104];
    tr.matrix_result[5].q[14] = mxu_if.mxu_lsu_int16_row5_data[119:112];
    tr.matrix_result[5].q[15] = mxu_if.mxu_lsu_int16_row5_data[127:120];
    tr.matrix_result[6].q[0] = mxu_if.mxu_lsu_int16_row6_data[7:0];
    tr.matrix_result[6].q[1] = mxu_if.mxu_lsu_int16_row6_data[15:8];
    tr.matrix_result[6].q[2] = mxu_if.mxu_lsu_int16_row6_data[23:16];
    tr.matrix_result[6].q[3] = mxu_if.mxu_lsu_int16_row6_data[31:24];
    tr.matrix_result[6].q[4] = mxu_if.mxu_lsu_int16_row6_data[39:32];
    tr.matrix_result[6].q[5] = mxu_if.mxu_lsu_int16_row6_data[47:40];
    tr.matrix_result[6].q[6] = mxu_if.mxu_lsu_int16_row6_data[55:48];
    tr.matrix_result[6].q[7] = mxu_if.mxu_lsu_int16_row6_data[63:56];
    tr.matrix_result[6].q[8] = mxu_if.mxu_lsu_int16_row6_data[71:64];
    tr.matrix_result[6].q[9] = mxu_if.mxu_lsu_int16_row6_data[79:72];
    tr.matrix_result[6].q[10] = mxu_if.mxu_lsu_int16_row6_data[87:80];
    tr.matrix_result[6].q[11] = mxu_if.mxu_lsu_int16_row6_data[95:88];
    tr.matrix_result[6].q[12] = mxu_if.mxu_lsu_int16_row6_data[103:96];
    tr.matrix_result[6].q[13] = mxu_if.mxu_lsu_int16_row6_data[111:104];
    tr.matrix_result[6].q[14] = mxu_if.mxu_lsu_int16_row6_data[119:112];
    tr.matrix_result[6].q[15] = mxu_if.mxu_lsu_int16_row6_data[127:120];
    tr.matrix_result[7].q[0] = mxu_if.mxu_lsu_int16_row7_data[7:0];
    tr.matrix_result[7].q[1] = mxu_if.mxu_lsu_int16_row7_data[15:8];
    tr.matrix_result[7].q[2] = mxu_if.mxu_lsu_int16_row7_data[23:16];
    tr.matrix_result[7].q[3] = mxu_if.mxu_lsu_int16_row7_data[31:24];
    tr.matrix_result[7].q[4] = mxu_if.mxu_lsu_int16_row7_data[39:32];
    tr.matrix_result[7].q[5] = mxu_if.mxu_lsu_int16_row7_data[47:40];
    tr.matrix_result[7].q[6] = mxu_if.mxu_lsu_int16_row7_data[55:48];
    tr.matrix_result[7].q[7] = mxu_if.mxu_lsu_int16_row7_data[63:56];
    tr.matrix_result[7].q[8] = mxu_if.mxu_lsu_int16_row7_data[71:64];
    tr.matrix_result[7].q[9] = mxu_if.mxu_lsu_int16_row7_data[79:72];
    tr.matrix_result[7].q[10] = mxu_if.mxu_lsu_int16_row7_data[87:80];
    tr.matrix_result[7].q[11] = mxu_if.mxu_lsu_int16_row7_data[95:88];
    tr.matrix_result[7].q[12] = mxu_if.mxu_lsu_int16_row7_data[103:96];
    tr.matrix_result[7].q[13] = mxu_if.mxu_lsu_int16_row7_data[111:104];
    tr.matrix_result[7].q[14] = mxu_if.mxu_lsu_int16_row7_data[119:112];
    tr.matrix_result[7].q[15] = mxu_if.mxu_lsu_int16_row7_data[127:120];
    tr.matrix_result[8].q[0] = mxu_if.mxu_lsu_int16_row8_data[7:0];
    tr.matrix_result[8].q[1] = mxu_if.mxu_lsu_int16_row8_data[15:8];
    tr.matrix_result[8].q[2] = mxu_if.mxu_lsu_int16_row8_data[23:16];
    tr.matrix_result[8].q[3] = mxu_if.mxu_lsu_int16_row8_data[31:24];
    tr.matrix_result[8].q[4] = mxu_if.mxu_lsu_int16_row8_data[39:32];
    tr.matrix_result[8].q[5] = mxu_if.mxu_lsu_int16_row8_data[47:40];
    tr.matrix_result[8].q[6] = mxu_if.mxu_lsu_int16_row8_data[55:48];
    tr.matrix_result[8].q[7] = mxu_if.mxu_lsu_int16_row8_data[63:56];
    tr.matrix_result[8].q[8] = mxu_if.mxu_lsu_int16_row8_data[71:64];
    tr.matrix_result[8].q[9] = mxu_if.mxu_lsu_int16_row8_data[79:72];
    tr.matrix_result[8].q[10] = mxu_if.mxu_lsu_int16_row8_data[87:80];
    tr.matrix_result[8].q[11] = mxu_if.mxu_lsu_int16_row8_data[95:88];
    tr.matrix_result[8].q[12] = mxu_if.mxu_lsu_int16_row8_data[103:96];
    tr.matrix_result[8].q[13] = mxu_if.mxu_lsu_int16_row8_data[111:104];
    tr.matrix_result[8].q[14] = mxu_if.mxu_lsu_int16_row8_data[119:112];
    tr.matrix_result[8].q[15] = mxu_if.mxu_lsu_int16_row8_data[127:120];
    tr.matrix_result[9].q[0] = mxu_if.mxu_lsu_int16_row9_data[7:0];
    tr.matrix_result[9].q[1] = mxu_if.mxu_lsu_int16_row9_data[15:8];
    tr.matrix_result[9].q[2] = mxu_if.mxu_lsu_int16_row9_data[23:16];
    tr.matrix_result[9].q[3] = mxu_if.mxu_lsu_int16_row9_data[31:24];
    tr.matrix_result[9].q[4] = mxu_if.mxu_lsu_int16_row9_data[39:32];
    tr.matrix_result[9].q[5] = mxu_if.mxu_lsu_int16_row9_data[47:40];
    tr.matrix_result[9].q[6] = mxu_if.mxu_lsu_int16_row9_data[55:48];
    tr.matrix_result[9].q[7] = mxu_if.mxu_lsu_int16_row9_data[63:56];
    tr.matrix_result[9].q[8] = mxu_if.mxu_lsu_int16_row9_data[71:64];
    tr.matrix_result[9].q[9] = mxu_if.mxu_lsu_int16_row9_data[79:72];
    tr.matrix_result[9].q[10] = mxu_if.mxu_lsu_int16_row9_data[87:80];
    tr.matrix_result[9].q[11] = mxu_if.mxu_lsu_int16_row9_data[95:88];
    tr.matrix_result[9].q[12] = mxu_if.mxu_lsu_int16_row9_data[103:96];
    tr.matrix_result[9].q[13] = mxu_if.mxu_lsu_int16_row9_data[111:104];
    tr.matrix_result[9].q[14] = mxu_if.mxu_lsu_int16_row9_data[119:112];
    tr.matrix_result[9].q[15] = mxu_if.mxu_lsu_int16_row9_data[127:120];
    tr.matrix_result[10].q[0] = mxu_if.mxu_lsu_int16_row10_data[7:0];
    tr.matrix_result[10].q[1] = mxu_if.mxu_lsu_int16_row10_data[15:8];
    tr.matrix_result[10].q[2] = mxu_if.mxu_lsu_int16_row10_data[23:16];
    tr.matrix_result[10].q[3] = mxu_if.mxu_lsu_int16_row10_data[31:24];
    tr.matrix_result[10].q[4] = mxu_if.mxu_lsu_int16_row10_data[39:32];
    tr.matrix_result[10].q[5] = mxu_if.mxu_lsu_int16_row10_data[47:40];
    tr.matrix_result[10].q[6] = mxu_if.mxu_lsu_int16_row10_data[55:48];
    tr.matrix_result[10].q[7] = mxu_if.mxu_lsu_int16_row10_data[63:56];
    tr.matrix_result[10].q[8] = mxu_if.mxu_lsu_int16_row10_data[71:64];
    tr.matrix_result[10].q[9] = mxu_if.mxu_lsu_int16_row10_data[79:72];
    tr.matrix_result[10].q[10] = mxu_if.mxu_lsu_int16_row10_data[87:80];
    tr.matrix_result[10].q[11] = mxu_if.mxu_lsu_int16_row10_data[95:88];
    tr.matrix_result[10].q[12] = mxu_if.mxu_lsu_int16_row10_data[103:96];
    tr.matrix_result[10].q[13] = mxu_if.mxu_lsu_int16_row10_data[111:104];
    tr.matrix_result[10].q[14] = mxu_if.mxu_lsu_int16_row10_data[119:112];
    tr.matrix_result[10].q[15] = mxu_if.mxu_lsu_int16_row10_data[127:120];
    tr.matrix_result[11].q[0] = mxu_if.mxu_lsu_int16_row11_data[7:0];
    tr.matrix_result[11].q[1] = mxu_if.mxu_lsu_int16_row11_data[15:8];
    tr.matrix_result[11].q[2] = mxu_if.mxu_lsu_int16_row11_data[23:16];
    tr.matrix_result[11].q[3] = mxu_if.mxu_lsu_int16_row11_data[31:24];
    tr.matrix_result[11].q[4] = mxu_if.mxu_lsu_int16_row11_data[39:32];
    tr.matrix_result[11].q[5] = mxu_if.mxu_lsu_int16_row11_data[47:40];
    tr.matrix_result[11].q[6] = mxu_if.mxu_lsu_int16_row11_data[55:48];
    tr.matrix_result[11].q[7] = mxu_if.mxu_lsu_int16_row11_data[63:56];
    tr.matrix_result[11].q[8] = mxu_if.mxu_lsu_int16_row11_data[71:64];
    tr.matrix_result[11].q[9] = mxu_if.mxu_lsu_int16_row11_data[79:72];
    tr.matrix_result[11].q[10] = mxu_if.mxu_lsu_int16_row11_data[87:80];
    tr.matrix_result[11].q[11] = mxu_if.mxu_lsu_int16_row11_data[95:88];
    tr.matrix_result[11].q[12] = mxu_if.mxu_lsu_int16_row11_data[103:96];
    tr.matrix_result[11].q[13] = mxu_if.mxu_lsu_int16_row11_data[111:104];
    tr.matrix_result[11].q[14] = mxu_if.mxu_lsu_int16_row11_data[119:112];
    tr.matrix_result[11].q[15] = mxu_if.mxu_lsu_int16_row11_data[127:120];
    tr.matrix_result[12].q[0] = mxu_if.mxu_lsu_int16_row12_data[7:0];
    tr.matrix_result[12].q[1] = mxu_if.mxu_lsu_int16_row12_data[15:8];
    tr.matrix_result[12].q[2] = mxu_if.mxu_lsu_int16_row12_data[23:16];
    tr.matrix_result[12].q[3] = mxu_if.mxu_lsu_int16_row12_data[31:24];
    tr.matrix_result[12].q[4] = mxu_if.mxu_lsu_int16_row12_data[39:32];
    tr.matrix_result[12].q[5] = mxu_if.mxu_lsu_int16_row12_data[47:40];
    tr.matrix_result[12].q[6] = mxu_if.mxu_lsu_int16_row12_data[55:48];
    tr.matrix_result[12].q[7] = mxu_if.mxu_lsu_int16_row12_data[63:56];
    tr.matrix_result[12].q[8] = mxu_if.mxu_lsu_int16_row12_data[71:64];
    tr.matrix_result[12].q[9] = mxu_if.mxu_lsu_int16_row12_data[79:72];
    tr.matrix_result[12].q[10] = mxu_if.mxu_lsu_int16_row12_data[87:80];
    tr.matrix_result[12].q[11] = mxu_if.mxu_lsu_int16_row12_data[95:88];
    tr.matrix_result[12].q[12] = mxu_if.mxu_lsu_int16_row12_data[103:96];
    tr.matrix_result[12].q[13] = mxu_if.mxu_lsu_int16_row12_data[111:104];
    tr.matrix_result[12].q[14] = mxu_if.mxu_lsu_int16_row12_data[119:112];
    tr.matrix_result[12].q[15] = mxu_if.mxu_lsu_int16_row12_data[127:120];
    tr.matrix_result[13].q[0] = mxu_if.mxu_lsu_int16_row13_data[7:0];
    tr.matrix_result[13].q[1] = mxu_if.mxu_lsu_int16_row13_data[15:8];
    tr.matrix_result[13].q[2] = mxu_if.mxu_lsu_int16_row13_data[23:16];
    tr.matrix_result[13].q[3] = mxu_if.mxu_lsu_int16_row13_data[31:24];
    tr.matrix_result[13].q[4] = mxu_if.mxu_lsu_int16_row13_data[39:32];
    tr.matrix_result[13].q[5] = mxu_if.mxu_lsu_int16_row13_data[47:40];
    tr.matrix_result[13].q[6] = mxu_if.mxu_lsu_int16_row13_data[55:48];
    tr.matrix_result[13].q[7] = mxu_if.mxu_lsu_int16_row13_data[63:56];
    tr.matrix_result[13].q[8] = mxu_if.mxu_lsu_int16_row13_data[71:64];
    tr.matrix_result[13].q[9] = mxu_if.mxu_lsu_int16_row13_data[79:72];
    tr.matrix_result[13].q[10] = mxu_if.mxu_lsu_int16_row13_data[87:80];
    tr.matrix_result[13].q[11] = mxu_if.mxu_lsu_int16_row13_data[95:88];
    tr.matrix_result[13].q[12] = mxu_if.mxu_lsu_int16_row13_data[103:96];
    tr.matrix_result[13].q[13] = mxu_if.mxu_lsu_int16_row13_data[111:104];
    tr.matrix_result[13].q[14] = mxu_if.mxu_lsu_int16_row13_data[119:112];
    tr.matrix_result[13].q[15] = mxu_if.mxu_lsu_int16_row13_data[127:120];
    tr.matrix_result[14].q[0] = mxu_if.mxu_lsu_int16_row14_data[7:0];
    tr.matrix_result[14].q[1] = mxu_if.mxu_lsu_int16_row14_data[15:8];
    tr.matrix_result[14].q[2] = mxu_if.mxu_lsu_int16_row14_data[23:16];
    tr.matrix_result[14].q[3] = mxu_if.mxu_lsu_int16_row14_data[31:24];
    tr.matrix_result[14].q[4] = mxu_if.mxu_lsu_int16_row14_data[39:32];
    tr.matrix_result[14].q[5] = mxu_if.mxu_lsu_int16_row14_data[47:40];
    tr.matrix_result[14].q[6] = mxu_if.mxu_lsu_int16_row14_data[55:48];
    tr.matrix_result[14].q[7] = mxu_if.mxu_lsu_int16_row14_data[63:56];
    tr.matrix_result[14].q[8] = mxu_if.mxu_lsu_int16_row14_data[71:64];
    tr.matrix_result[14].q[9] = mxu_if.mxu_lsu_int16_row14_data[79:72];
    tr.matrix_result[14].q[10] = mxu_if.mxu_lsu_int16_row14_data[87:80];
    tr.matrix_result[14].q[11] = mxu_if.mxu_lsu_int16_row14_data[95:88];
    tr.matrix_result[14].q[12] = mxu_if.mxu_lsu_int16_row14_data[103:96];
    tr.matrix_result[14].q[13] = mxu_if.mxu_lsu_int16_row14_data[111:104];
    tr.matrix_result[14].q[14] = mxu_if.mxu_lsu_int16_row14_data[119:112];
    tr.matrix_result[14].q[15] = mxu_if.mxu_lsu_int16_row14_data[127:120];
    tr.matrix_result[15].q[0] = mxu_if.mxu_lsu_int16_row15_data[7:0];
    tr.matrix_result[15].q[1] = mxu_if.mxu_lsu_int16_row15_data[15:8];
    tr.matrix_result[15].q[2] = mxu_if.mxu_lsu_int16_row15_data[23:16];
    tr.matrix_result[15].q[3] = mxu_if.mxu_lsu_int16_row15_data[31:24];
    tr.matrix_result[15].q[4] = mxu_if.mxu_lsu_int16_row15_data[39:32];
    tr.matrix_result[15].q[5] = mxu_if.mxu_lsu_int16_row15_data[47:40];
    tr.matrix_result[15].q[6] = mxu_if.mxu_lsu_int16_row15_data[55:48];
    tr.matrix_result[15].q[7] = mxu_if.mxu_lsu_int16_row15_data[63:56];
    tr.matrix_result[15].q[8] = mxu_if.mxu_lsu_int16_row15_data[71:64];
    tr.matrix_result[15].q[9] = mxu_if.mxu_lsu_int16_row15_data[79:72];
    tr.matrix_result[15].q[10] = mxu_if.mxu_lsu_int16_row15_data[87:80];
    tr.matrix_result[15].q[11] = mxu_if.mxu_lsu_int16_row15_data[95:88];
    tr.matrix_result[15].q[12] = mxu_if.mxu_lsu_int16_row15_data[103:96];
    tr.matrix_result[15].q[13] = mxu_if.mxu_lsu_int16_row15_data[111:104];
    tr.matrix_result[15].q[14] = mxu_if.mxu_lsu_int16_row15_data[119:112];
    tr.matrix_result[15].q[15] = mxu_if.mxu_lsu_int16_row15_data[127:120];

endtask
