interface axi_wr_intf(
);

endinterface