class mxu_output_monitor extends uvm_monitor;

    virtual mxu_intf mxu_if;
    uvm_analysis_port #(mxu_tr) ap;

    `uvm_component_utils(mxu_output_monitor)
    function new(string name = "mxu_output_monitor", uvm_component parent = null);
       super.new(name, parent);
    endfunction //new()
    
    extern virtual task build_phase(uvm_phase phase);
    extern virtual task main_phase(uvm_phase phase);
    
    extern virtual task collect_matrix_out(mxu_tr tr);

endclass //mxu_output_monitor extends superClass

task mxu_output_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual mxu_intf)::get(this, "", "mxu_if", mxu_if))begin
        `uvm_fatal("mxu_output_monitor", "mxu output_monitor fail to get mxu if")
    end
    ap = new("ap", this);
endtask

task mxu_output_monitor::main_phase(uvm_phase phase);
    mxu_tr tr;

    tr = new("tr");

    while (1) begin 
        this.collect_matrix(tr);
        ap.write(tr);
    end

endtask

task mxu_output_monitor::collect_matrix_out(mxu_tr tr);

    while(1)begin
        @(posedge mxu_if.clk);
        if(mxu_if.lsu_mxu_vld) break;
    end

    tr.clear_result();
    @(posedge mxu_if.clk);
    wait(mxu_if.mxu_lsu_data_rdy) 
    tr.matrix_result[0][0] = mxu_if.mxu_lsu_int16_row0_data[7:0];
    tr.matrix_result[0][1] = mxu_if.mxu_lsu_int16_row0_data[15:8];
    tr.matrix_result[0][2] = mxu_if.mxu_lsu_int16_row0_data[23:16];
    tr.matrix_result[0][3] = mxu_if.mxu_lsu_int16_row0_data[31:24];
    tr.matrix_result[0][4] = mxu_if.mxu_lsu_int16_row0_data[39:32];
    tr.matrix_result[0][5] = mxu_if.mxu_lsu_int16_row0_data[47:40];
    tr.matrix_result[0][6] = mxu_if.mxu_lsu_int16_row0_data[55:48];
    tr.matrix_result[0][7] = mxu_if.mxu_lsu_int16_row0_data[63:56];
    tr.matrix_result[0][8] = mxu_if.mxu_lsu_int16_row0_data[71:64];
    tr.matrix_result[0][9] = mxu_if.mxu_lsu_int16_row0_data[79:72];
    tr.matrix_result[0][10] = mxu_if.mxu_lsu_int16_row0_data[87:80];
    tr.matrix_result[0][11] = mxu_if.mxu_lsu_int16_row0_data[95:88];
    tr.matrix_result[0][12] = mxu_if.mxu_lsu_int16_row0_data[103:96];
    tr.matrix_result[0][13] = mxu_if.mxu_lsu_int16_row0_data[111:104];
    tr.matrix_result[0][14] = mxu_if.mxu_lsu_int16_row0_data[119:112];
    tr.matrix_result[0][15] = mxu_if.mxu_lsu_int16_row0_data[127:120];
    tr.matrix_result[1][0] = mxu_if.mxu_lsu_int16_row1_data[7:0];
    tr.matrix_result[1][1] = mxu_if.mxu_lsu_int16_row1_data[15:8];
    tr.matrix_result[1][2] = mxu_if.mxu_lsu_int16_row1_data[23:16];
    tr.matrix_result[1][3] = mxu_if.mxu_lsu_int16_row1_data[31:24];
    tr.matrix_result[1][4] = mxu_if.mxu_lsu_int16_row1_data[39:32];
    tr.matrix_result[1][5] = mxu_if.mxu_lsu_int16_row1_data[47:40];
    tr.matrix_result[1][6] = mxu_if.mxu_lsu_int16_row1_data[55:48];
    tr.matrix_result[1][7] = mxu_if.mxu_lsu_int16_row1_data[63:56];
    tr.matrix_result[1][8] = mxu_if.mxu_lsu_int16_row1_data[71:64];
    tr.matrix_result[1][9] = mxu_if.mxu_lsu_int16_row1_data[79:72];
    tr.matrix_result[1][10] = mxu_if.mxu_lsu_int16_row1_data[87:80];
    tr.matrix_result[1][11] = mxu_if.mxu_lsu_int16_row1_data[95:88];
    tr.matrix_result[1][12] = mxu_if.mxu_lsu_int16_row1_data[103:96];
    tr.matrix_result[1][13] = mxu_if.mxu_lsu_int16_row1_data[111:104];
    tr.matrix_result[1][14] = mxu_if.mxu_lsu_int16_row1_data[119:112];
    tr.matrix_result[1][15] = mxu_if.mxu_lsu_int16_row1_data[127:120];
    tr.matrix_result[2][0] = mxu_if.mxu_lsu_int16_row2_data[7:0];
    tr.matrix_result[2][1] = mxu_if.mxu_lsu_int16_row2_data[15:8];
    tr.matrix_result[2][2] = mxu_if.mxu_lsu_int16_row2_data[23:16];
    tr.matrix_result[2][3] = mxu_if.mxu_lsu_int16_row2_data[31:24];
    tr.matrix_result[2][4] = mxu_if.mxu_lsu_int16_row2_data[39:32];
    tr.matrix_result[2][5] = mxu_if.mxu_lsu_int16_row2_data[47:40];
    tr.matrix_result[2][6] = mxu_if.mxu_lsu_int16_row2_data[55:48];
    tr.matrix_result[2][7] = mxu_if.mxu_lsu_int16_row2_data[63:56];
    tr.matrix_result[2][8] = mxu_if.mxu_lsu_int16_row2_data[71:64];
    tr.matrix_result[2][9] = mxu_if.mxu_lsu_int16_row2_data[79:72];
    tr.matrix_result[2][10] = mxu_if.mxu_lsu_int16_row2_data[87:80];
    tr.matrix_result[2][11] = mxu_if.mxu_lsu_int16_row2_data[95:88];
    tr.matrix_result[2][12] = mxu_if.mxu_lsu_int16_row2_data[103:96];
    tr.matrix_result[2][13] = mxu_if.mxu_lsu_int16_row2_data[111:104];
    tr.matrix_result[2][14] = mxu_if.mxu_lsu_int16_row2_data[119:112];
    tr.matrix_result[2][15] = mxu_if.mxu_lsu_int16_row2_data[127:120];
    tr.matrix_result[3][0] = mxu_if.mxu_lsu_int16_row3_data[7:0];
    tr.matrix_result[3][1] = mxu_if.mxu_lsu_int16_row3_data[15:8];
    tr.matrix_result[3][2] = mxu_if.mxu_lsu_int16_row3_data[23:16];
    tr.matrix_result[3][3] = mxu_if.mxu_lsu_int16_row3_data[31:24];
    tr.matrix_result[3][4] = mxu_if.mxu_lsu_int16_row3_data[39:32];
    tr.matrix_result[3][5] = mxu_if.mxu_lsu_int16_row3_data[47:40];
    tr.matrix_result[3][6] = mxu_if.mxu_lsu_int16_row3_data[55:48];
    tr.matrix_result[3][7] = mxu_if.mxu_lsu_int16_row3_data[63:56];
    tr.matrix_result[3][8] = mxu_if.mxu_lsu_int16_row3_data[71:64];
    tr.matrix_result[3][9] = mxu_if.mxu_lsu_int16_row3_data[79:72];
    tr.matrix_result[3][10] = mxu_if.mxu_lsu_int16_row3_data[87:80];
    tr.matrix_result[3][11] = mxu_if.mxu_lsu_int16_row3_data[95:88];
    tr.matrix_result[3][12] = mxu_if.mxu_lsu_int16_row3_data[103:96];
    tr.matrix_result[3][13] = mxu_if.mxu_lsu_int16_row3_data[111:104];
    tr.matrix_result[3][14] = mxu_if.mxu_lsu_int16_row3_data[119:112];
    tr.matrix_result[3][15] = mxu_if.mxu_lsu_int16_row3_data[127:120];
    tr.matrix_result[4][0] = mxu_if.mxu_lsu_int16_row4_data[7:0];
    tr.matrix_result[4][1] = mxu_if.mxu_lsu_int16_row4_data[15:8];
    tr.matrix_result[4][2] = mxu_if.mxu_lsu_int16_row4_data[23:16];
    tr.matrix_result[4][3] = mxu_if.mxu_lsu_int16_row4_data[31:24];
    tr.matrix_result[4][4] = mxu_if.mxu_lsu_int16_row4_data[39:32];
    tr.matrix_result[4][5] = mxu_if.mxu_lsu_int16_row4_data[47:40];
    tr.matrix_result[4][6] = mxu_if.mxu_lsu_int16_row4_data[55:48];
    tr.matrix_result[4][7] = mxu_if.mxu_lsu_int16_row4_data[63:56];
    tr.matrix_result[4][8] = mxu_if.mxu_lsu_int16_row4_data[71:64];
    tr.matrix_result[4][9] = mxu_if.mxu_lsu_int16_row4_data[79:72];
    tr.matrix_result[4][10] = mxu_if.mxu_lsu_int16_row4_data[87:80];
    tr.matrix_result[4][11] = mxu_if.mxu_lsu_int16_row4_data[95:88];
    tr.matrix_result[4][12] = mxu_if.mxu_lsu_int16_row4_data[103:96];
    tr.matrix_result[4][13] = mxu_if.mxu_lsu_int16_row4_data[111:104];
    tr.matrix_result[4][14] = mxu_if.mxu_lsu_int16_row4_data[119:112];
    tr.matrix_result[4][15] = mxu_if.mxu_lsu_int16_row4_data[127:120];
    tr.matrix_result[5][0] = mxu_if.mxu_lsu_int16_row5_data[7:0];
    tr.matrix_result[5][1] = mxu_if.mxu_lsu_int16_row5_data[15:8];
    tr.matrix_result[5][2] = mxu_if.mxu_lsu_int16_row5_data[23:16];
    tr.matrix_result[5][3] = mxu_if.mxu_lsu_int16_row5_data[31:24];
    tr.matrix_result[5][4] = mxu_if.mxu_lsu_int16_row5_data[39:32];
    tr.matrix_result[5][5] = mxu_if.mxu_lsu_int16_row5_data[47:40];
    tr.matrix_result[5][6] = mxu_if.mxu_lsu_int16_row5_data[55:48];
    tr.matrix_result[5][7] = mxu_if.mxu_lsu_int16_row5_data[63:56];
    tr.matrix_result[5][8] = mxu_if.mxu_lsu_int16_row5_data[71:64];
    tr.matrix_result[5][9] = mxu_if.mxu_lsu_int16_row5_data[79:72];
    tr.matrix_result[5][10] = mxu_if.mxu_lsu_int16_row5_data[87:80];
    tr.matrix_result[5][11] = mxu_if.mxu_lsu_int16_row5_data[95:88];
    tr.matrix_result[5][12] = mxu_if.mxu_lsu_int16_row5_data[103:96];
    tr.matrix_result[5][13] = mxu_if.mxu_lsu_int16_row5_data[111:104];
    tr.matrix_result[5][14] = mxu_if.mxu_lsu_int16_row5_data[119:112];
    tr.matrix_result[5][15] = mxu_if.mxu_lsu_int16_row5_data[127:120];
    tr.matrix_result[6][0] = mxu_if.mxu_lsu_int16_row6_data[7:0];
    tr.matrix_result[6][1] = mxu_if.mxu_lsu_int16_row6_data[15:8];
    tr.matrix_result[6][2] = mxu_if.mxu_lsu_int16_row6_data[23:16];
    tr.matrix_result[6][3] = mxu_if.mxu_lsu_int16_row6_data[31:24];
    tr.matrix_result[6][4] = mxu_if.mxu_lsu_int16_row6_data[39:32];
    tr.matrix_result[6][5] = mxu_if.mxu_lsu_int16_row6_data[47:40];
    tr.matrix_result[6][6] = mxu_if.mxu_lsu_int16_row6_data[55:48];
    tr.matrix_result[6][7] = mxu_if.mxu_lsu_int16_row6_data[63:56];
    tr.matrix_result[6][8] = mxu_if.mxu_lsu_int16_row6_data[71:64];
    tr.matrix_result[6][9] = mxu_if.mxu_lsu_int16_row6_data[79:72];
    tr.matrix_result[6][10] = mxu_if.mxu_lsu_int16_row6_data[87:80];
    tr.matrix_result[6][11] = mxu_if.mxu_lsu_int16_row6_data[95:88];
    tr.matrix_result[6][12] = mxu_if.mxu_lsu_int16_row6_data[103:96];
    tr.matrix_result[6][13] = mxu_if.mxu_lsu_int16_row6_data[111:104];
    tr.matrix_result[6][14] = mxu_if.mxu_lsu_int16_row6_data[119:112];
    tr.matrix_result[6][15] = mxu_if.mxu_lsu_int16_row6_data[127:120];
    tr.matrix_result[7][0] = mxu_if.mxu_lsu_int16_row7_data[7:0];
    tr.matrix_result[7][1] = mxu_if.mxu_lsu_int16_row7_data[15:8];
    tr.matrix_result[7][2] = mxu_if.mxu_lsu_int16_row7_data[23:16];
    tr.matrix_result[7][3] = mxu_if.mxu_lsu_int16_row7_data[31:24];
    tr.matrix_result[7][4] = mxu_if.mxu_lsu_int16_row7_data[39:32];
    tr.matrix_result[7][5] = mxu_if.mxu_lsu_int16_row7_data[47:40];
    tr.matrix_result[7][6] = mxu_if.mxu_lsu_int16_row7_data[55:48];
    tr.matrix_result[7][7] = mxu_if.mxu_lsu_int16_row7_data[63:56];
    tr.matrix_result[7][8] = mxu_if.mxu_lsu_int16_row7_data[71:64];
    tr.matrix_result[7][9] = mxu_if.mxu_lsu_int16_row7_data[79:72];
    tr.matrix_result[7][10] = mxu_if.mxu_lsu_int16_row7_data[87:80];
    tr.matrix_result[7][11] = mxu_if.mxu_lsu_int16_row7_data[95:88];
    tr.matrix_result[7][12] = mxu_if.mxu_lsu_int16_row7_data[103:96];
    tr.matrix_result[7][13] = mxu_if.mxu_lsu_int16_row7_data[111:104];
    tr.matrix_result[7][14] = mxu_if.mxu_lsu_int16_row7_data[119:112];
    tr.matrix_result[7][15] = mxu_if.mxu_lsu_int16_row7_data[127:120];
    tr.matrix_result[8][0] = mxu_if.mxu_lsu_int16_row8_data[7:0];
    tr.matrix_result[8][1] = mxu_if.mxu_lsu_int16_row8_data[15:8];
    tr.matrix_result[8][2] = mxu_if.mxu_lsu_int16_row8_data[23:16];
    tr.matrix_result[8][3] = mxu_if.mxu_lsu_int16_row8_data[31:24];
    tr.matrix_result[8][4] = mxu_if.mxu_lsu_int16_row8_data[39:32];
    tr.matrix_result[8][5] = mxu_if.mxu_lsu_int16_row8_data[47:40];
    tr.matrix_result[8][6] = mxu_if.mxu_lsu_int16_row8_data[55:48];
    tr.matrix_result[8][7] = mxu_if.mxu_lsu_int16_row8_data[63:56];
    tr.matrix_result[8][8] = mxu_if.mxu_lsu_int16_row8_data[71:64];
    tr.matrix_result[8][9] = mxu_if.mxu_lsu_int16_row8_data[79:72];
    tr.matrix_result[8][10] = mxu_if.mxu_lsu_int16_row8_data[87:80];
    tr.matrix_result[8][11] = mxu_if.mxu_lsu_int16_row8_data[95:88];
    tr.matrix_result[8][12] = mxu_if.mxu_lsu_int16_row8_data[103:96];
    tr.matrix_result[8][13] = mxu_if.mxu_lsu_int16_row8_data[111:104];
    tr.matrix_result[8][14] = mxu_if.mxu_lsu_int16_row8_data[119:112];
    tr.matrix_result[8][15] = mxu_if.mxu_lsu_int16_row8_data[127:120];
    tr.matrix_result[9][0] = mxu_if.mxu_lsu_int16_row9_data[7:0];
    tr.matrix_result[9][1] = mxu_if.mxu_lsu_int16_row9_data[15:8];
    tr.matrix_result[9][2] = mxu_if.mxu_lsu_int16_row9_data[23:16];
    tr.matrix_result[9][3] = mxu_if.mxu_lsu_int16_row9_data[31:24];
    tr.matrix_result[9][4] = mxu_if.mxu_lsu_int16_row9_data[39:32];
    tr.matrix_result[9][5] = mxu_if.mxu_lsu_int16_row9_data[47:40];
    tr.matrix_result[9][6] = mxu_if.mxu_lsu_int16_row9_data[55:48];
    tr.matrix_result[9][7] = mxu_if.mxu_lsu_int16_row9_data[63:56];
    tr.matrix_result[9][8] = mxu_if.mxu_lsu_int16_row9_data[71:64];
    tr.matrix_result[9][9] = mxu_if.mxu_lsu_int16_row9_data[79:72];
    tr.matrix_result[9][10] = mxu_if.mxu_lsu_int16_row9_data[87:80];
    tr.matrix_result[9][11] = mxu_if.mxu_lsu_int16_row9_data[95:88];
    tr.matrix_result[9][12] = mxu_if.mxu_lsu_int16_row9_data[103:96];
    tr.matrix_result[9][13] = mxu_if.mxu_lsu_int16_row9_data[111:104];
    tr.matrix_result[9][14] = mxu_if.mxu_lsu_int16_row9_data[119:112];
    tr.matrix_result[9][15] = mxu_if.mxu_lsu_int16_row9_data[127:120];
    tr.matrix_result[10][0] = mxu_if.mxu_lsu_int16_row10_data[7:0];
    tr.matrix_result[10][1] = mxu_if.mxu_lsu_int16_row10_data[15:8];
    tr.matrix_result[10][2] = mxu_if.mxu_lsu_int16_row10_data[23:16];
    tr.matrix_result[10][3] = mxu_if.mxu_lsu_int16_row10_data[31:24];
    tr.matrix_result[10][4] = mxu_if.mxu_lsu_int16_row10_data[39:32];
    tr.matrix_result[10][5] = mxu_if.mxu_lsu_int16_row10_data[47:40];
    tr.matrix_result[10][6] = mxu_if.mxu_lsu_int16_row10_data[55:48];
    tr.matrix_result[10][7] = mxu_if.mxu_lsu_int16_row10_data[63:56];
    tr.matrix_result[10][8] = mxu_if.mxu_lsu_int16_row10_data[71:64];
    tr.matrix_result[10][9] = mxu_if.mxu_lsu_int16_row10_data[79:72];
    tr.matrix_result[10][10] = mxu_if.mxu_lsu_int16_row10_data[87:80];
    tr.matrix_result[10][11] = mxu_if.mxu_lsu_int16_row10_data[95:88];
    tr.matrix_result[10][12] = mxu_if.mxu_lsu_int16_row10_data[103:96];
    tr.matrix_result[10][13] = mxu_if.mxu_lsu_int16_row10_data[111:104];
    tr.matrix_result[10][14] = mxu_if.mxu_lsu_int16_row10_data[119:112];
    tr.matrix_result[10][15] = mxu_if.mxu_lsu_int16_row10_data[127:120];
    tr.matrix_result[11][0] = mxu_if.mxu_lsu_int16_row11_data[7:0];
    tr.matrix_result[11][1] = mxu_if.mxu_lsu_int16_row11_data[15:8];
    tr.matrix_result[11][2] = mxu_if.mxu_lsu_int16_row11_data[23:16];
    tr.matrix_result[11][3] = mxu_if.mxu_lsu_int16_row11_data[31:24];
    tr.matrix_result[11][4] = mxu_if.mxu_lsu_int16_row11_data[39:32];
    tr.matrix_result[11][5] = mxu_if.mxu_lsu_int16_row11_data[47:40];
    tr.matrix_result[11][6] = mxu_if.mxu_lsu_int16_row11_data[55:48];
    tr.matrix_result[11][7] = mxu_if.mxu_lsu_int16_row11_data[63:56];
    tr.matrix_result[11][8] = mxu_if.mxu_lsu_int16_row11_data[71:64];
    tr.matrix_result[11][9] = mxu_if.mxu_lsu_int16_row11_data[79:72];
    tr.matrix_result[11][10] = mxu_if.mxu_lsu_int16_row11_data[87:80];
    tr.matrix_result[11][11] = mxu_if.mxu_lsu_int16_row11_data[95:88];
    tr.matrix_result[11][12] = mxu_if.mxu_lsu_int16_row11_data[103:96];
    tr.matrix_result[11][13] = mxu_if.mxu_lsu_int16_row11_data[111:104];
    tr.matrix_result[11][14] = mxu_if.mxu_lsu_int16_row11_data[119:112];
    tr.matrix_result[11][15] = mxu_if.mxu_lsu_int16_row11_data[127:120];
    tr.matrix_result[12][0] = mxu_if.mxu_lsu_int16_row12_data[7:0];
    tr.matrix_result[12][1] = mxu_if.mxu_lsu_int16_row12_data[15:8];
    tr.matrix_result[12][2] = mxu_if.mxu_lsu_int16_row12_data[23:16];
    tr.matrix_result[12][3] = mxu_if.mxu_lsu_int16_row12_data[31:24];
    tr.matrix_result[12][4] = mxu_if.mxu_lsu_int16_row12_data[39:32];
    tr.matrix_result[12][5] = mxu_if.mxu_lsu_int16_row12_data[47:40];
    tr.matrix_result[12][6] = mxu_if.mxu_lsu_int16_row12_data[55:48];
    tr.matrix_result[12][7] = mxu_if.mxu_lsu_int16_row12_data[63:56];
    tr.matrix_result[12][8] = mxu_if.mxu_lsu_int16_row12_data[71:64];
    tr.matrix_result[12][9] = mxu_if.mxu_lsu_int16_row12_data[79:72];
    tr.matrix_result[12][10] = mxu_if.mxu_lsu_int16_row12_data[87:80];
    tr.matrix_result[12][11] = mxu_if.mxu_lsu_int16_row12_data[95:88];
    tr.matrix_result[12][12] = mxu_if.mxu_lsu_int16_row12_data[103:96];
    tr.matrix_result[12][13] = mxu_if.mxu_lsu_int16_row12_data[111:104];
    tr.matrix_result[12][14] = mxu_if.mxu_lsu_int16_row12_data[119:112];
    tr.matrix_result[12][15] = mxu_if.mxu_lsu_int16_row12_data[127:120];
    tr.matrix_result[13][0] = mxu_if.mxu_lsu_int16_row13_data[7:0];
    tr.matrix_result[13][1] = mxu_if.mxu_lsu_int16_row13_data[15:8];
    tr.matrix_result[13][2] = mxu_if.mxu_lsu_int16_row13_data[23:16];
    tr.matrix_result[13][3] = mxu_if.mxu_lsu_int16_row13_data[31:24];
    tr.matrix_result[13][4] = mxu_if.mxu_lsu_int16_row13_data[39:32];
    tr.matrix_result[13][5] = mxu_if.mxu_lsu_int16_row13_data[47:40];
    tr.matrix_result[13][6] = mxu_if.mxu_lsu_int16_row13_data[55:48];
    tr.matrix_result[13][7] = mxu_if.mxu_lsu_int16_row13_data[63:56];
    tr.matrix_result[13][8] = mxu_if.mxu_lsu_int16_row13_data[71:64];
    tr.matrix_result[13][9] = mxu_if.mxu_lsu_int16_row13_data[79:72];
    tr.matrix_result[13][10] = mxu_if.mxu_lsu_int16_row13_data[87:80];
    tr.matrix_result[13][11] = mxu_if.mxu_lsu_int16_row13_data[95:88];
    tr.matrix_result[13][12] = mxu_if.mxu_lsu_int16_row13_data[103:96];
    tr.matrix_result[13][13] = mxu_if.mxu_lsu_int16_row13_data[111:104];
    tr.matrix_result[13][14] = mxu_if.mxu_lsu_int16_row13_data[119:112];
    tr.matrix_result[13][15] = mxu_if.mxu_lsu_int16_row13_data[127:120];
    tr.matrix_result[14][0] = mxu_if.mxu_lsu_int16_row14_data[7:0];
    tr.matrix_result[14][1] = mxu_if.mxu_lsu_int16_row14_data[15:8];
    tr.matrix_result[14][2] = mxu_if.mxu_lsu_int16_row14_data[23:16];
    tr.matrix_result[14][3] = mxu_if.mxu_lsu_int16_row14_data[31:24];
    tr.matrix_result[14][4] = mxu_if.mxu_lsu_int16_row14_data[39:32];
    tr.matrix_result[14][5] = mxu_if.mxu_lsu_int16_row14_data[47:40];
    tr.matrix_result[14][6] = mxu_if.mxu_lsu_int16_row14_data[55:48];
    tr.matrix_result[14][7] = mxu_if.mxu_lsu_int16_row14_data[63:56];
    tr.matrix_result[14][8] = mxu_if.mxu_lsu_int16_row14_data[71:64];
    tr.matrix_result[14][9] = mxu_if.mxu_lsu_int16_row14_data[79:72];
    tr.matrix_result[14][10] = mxu_if.mxu_lsu_int16_row14_data[87:80];
    tr.matrix_result[14][11] = mxu_if.mxu_lsu_int16_row14_data[95:88];
    tr.matrix_result[14][12] = mxu_if.mxu_lsu_int16_row14_data[103:96];
    tr.matrix_result[14][13] = mxu_if.mxu_lsu_int16_row14_data[111:104];
    tr.matrix_result[14][14] = mxu_if.mxu_lsu_int16_row14_data[119:112];
    tr.matrix_result[14][15] = mxu_if.mxu_lsu_int16_row14_data[127:120];
    tr.matrix_result[15][0] = mxu_if.mxu_lsu_int16_row15_data[7:0];
    tr.matrix_result[15][1] = mxu_if.mxu_lsu_int16_row15_data[15:8];
    tr.matrix_result[15][2] = mxu_if.mxu_lsu_int16_row15_data[23:16];
    tr.matrix_result[15][3] = mxu_if.mxu_lsu_int16_row15_data[31:24];
    tr.matrix_result[15][4] = mxu_if.mxu_lsu_int16_row15_data[39:32];
    tr.matrix_result[15][5] = mxu_if.mxu_lsu_int16_row15_data[47:40];
    tr.matrix_result[15][6] = mxu_if.mxu_lsu_int16_row15_data[55:48];
    tr.matrix_result[15][7] = mxu_if.mxu_lsu_int16_row15_data[63:56];
    tr.matrix_result[15][8] = mxu_if.mxu_lsu_int16_row15_data[71:64];
    tr.matrix_result[15][9] = mxu_if.mxu_lsu_int16_row15_data[79:72];
    tr.matrix_result[15][10] = mxu_if.mxu_lsu_int16_row15_data[87:80];
    tr.matrix_result[15][11] = mxu_if.mxu_lsu_int16_row15_data[95:88];
    tr.matrix_result[15][12] = mxu_if.mxu_lsu_int16_row15_data[103:96];
    tr.matrix_result[15][13] = mxu_if.mxu_lsu_int16_row15_data[111:104];
    tr.matrix_result[15][14] = mxu_if.mxu_lsu_int16_row15_data[119:112];
    tr.matrix_result[15][15] = mxu_if.mxu_lsu_int16_row15_data[127:120];

endtask
