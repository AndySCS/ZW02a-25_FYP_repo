module act_mod(
    clk,
    rst_n,
    act_type,
    act_vld,
    row0_data,
    act_row0_vld,
    act_row0_data,
    row1_data,
    act_row1_vld,
    act_row1_data,
    row2_data,
    act_row2_vld,
    act_row2_data,
    row3_data,
    act_row3_vld,
    act_row3_data,
    row4_data,
    act_row4_vld,
    act_row4_data,
    row5_data,
    act_row5_vld,
    act_row5_data,
    row6_data,
    act_row6_vld,
    act_row6_data,
    row7_data,
    act_row7_vld,
    act_row7_data,
    row8_data,
    act_row8_vld,
    act_row8_data,
    row9_data,
    act_row9_vld,
    act_row9_data,
    row10_data,
    act_row10_vld,
    act_row10_data,
    row11_data,
    act_row11_vld,
    act_row11_data,
    row12_data,
    act_row12_vld,
    act_row12_data,
    row13_data,
    act_row13_vld,
    act_row13_data,
    row14_data,
    act_row14_vld,
    act_row14_data,
    row15_data,
    act_row15_vld,
    act_row15_data,
    act_busy
);
     
    input clk;
    input rst_n;
    input [1:0] act_type;
    input act_vld;
    input [255:0] row0_data;
    output [15:0] act_row0_vld;
    output [255:0] act_row0_data;
    input [255:0] row1_data;
    output [15:0] act_row1_vld;
    output [255:0] act_row1_data;
    input [255:0] row2_data;
    output [15:0] act_row2_vld;
    output [255:0] act_row2_data;
    input [255:0] row3_data;
    output [15:0] act_row3_vld;
    output [255:0] act_row3_data;
    input [255:0] row4_data;
    output [15:0] act_row4_vld;
    output [255:0] act_row4_data;
    input [255:0] row5_data;
    output [15:0] act_row5_vld;
    output [255:0] act_row5_data;
    input [255:0] row6_data;
    output [15:0] act_row6_vld;
    output [255:0] act_row6_data;
    input [255:0] row7_data;
    output [15:0] act_row7_vld;
    output [255:0] act_row7_data;
    input [255:0] row8_data;
    output [15:0] act_row8_vld;
    output [255:0] act_row8_data;
    input [255:0] row9_data;
    output [15:0] act_row9_vld;
    output [255:0] act_row9_data;
    input [255:0] row10_data;
    output [15:0] act_row10_vld;
    output [255:0] act_row10_data;
    input [255:0] row11_data;
    output [15:0] act_row11_vld;
    output [255:0] act_row11_data;
    input [255:0] row12_data;
    output [15:0] act_row12_vld;
    output [255:0] act_row12_data;
    input [255:0] row13_data;
    output [15:0] act_row13_vld;
    output [255:0] act_row13_data;
    input [255:0] row14_data;
    output [15:0] act_row14_vld;
    output [255:0] act_row14_data;
    input [255:0] row15_data;
    output [15:0] act_row15_vld;
    output [255:0] act_row15_data;
    output act_busy;

    assign act_busy = act_vld;

    assign act_row0_vld = {16{act_vld}};

    assign act_row0_data[15:0] = row0_data[15] ? 16'b0 : row0_data[15:0];
    assign act_row0_data[31:16] = row0_data[31] ? 16'b0 : row0_data[31:16];
    assign act_row0_data[47:32] = row0_data[47] ? 16'b0 : row0_data[47:32];
    assign act_row0_data[63:48] = row0_data[63] ? 16'b0 : row0_data[63:48];
    assign act_row0_data[79:64] = row0_data[79] ? 16'b0 : row0_data[79:64];
    assign act_row0_data[95:80] = row0_data[95] ? 16'b0 : row0_data[95:80];
    assign act_row0_data[111:96] = row0_data[111] ? 16'b0 : row0_data[111:96];
    assign act_row0_data[127:112] = row0_data[127] ? 16'b0 : row0_data[127:112];
    assign act_row0_data[143:128] = row0_data[143] ? 16'b0 : row0_data[143:128];
    assign act_row0_data[159:144] = row0_data[159] ? 16'b0 : row0_data[159:144];
    assign act_row0_data[175:160] = row0_data[175] ? 16'b0 : row0_data[175:160];
    assign act_row0_data[191:176] = row0_data[191] ? 16'b0 : row0_data[191:176];
    assign act_row0_data[207:192] = row0_data[207] ? 16'b0 : row0_data[207:192];
    assign act_row0_data[223:208] = row0_data[223] ? 16'b0 : row0_data[223:208];
    assign act_row0_data[239:224] = row0_data[239] ? 16'b0 : row0_data[239:224];
    assign act_row0_data[255:240] = row0_data[255] ? 16'b0 : row0_data[255:240];

    assign act_row1_vld = {16{act_vld}};

    assign act_row1_data[15:0] = row1_data[15] ? 16'b0 : row1_data[15:0];
    assign act_row1_data[31:16] = row1_data[31] ? 16'b0 : row1_data[31:16];
    assign act_row1_data[47:32] = row1_data[47] ? 16'b0 : row1_data[47:32];
    assign act_row1_data[63:48] = row1_data[63] ? 16'b0 : row1_data[63:48];
    assign act_row1_data[79:64] = row1_data[79] ? 16'b0 : row1_data[79:64];
    assign act_row1_data[95:80] = row1_data[95] ? 16'b0 : row1_data[95:80];
    assign act_row1_data[111:96] = row1_data[111] ? 16'b0 : row1_data[111:96];
    assign act_row1_data[127:112] = row1_data[127] ? 16'b0 : row1_data[127:112];
    assign act_row1_data[143:128] = row1_data[143] ? 16'b0 : row1_data[143:128];
    assign act_row1_data[159:144] = row1_data[159] ? 16'b0 : row1_data[159:144];
    assign act_row1_data[175:160] = row1_data[175] ? 16'b0 : row1_data[175:160];
    assign act_row1_data[191:176] = row1_data[191] ? 16'b0 : row1_data[191:176];
    assign act_row1_data[207:192] = row1_data[207] ? 16'b0 : row1_data[207:192];
    assign act_row1_data[223:208] = row1_data[223] ? 16'b0 : row1_data[223:208];
    assign act_row1_data[239:224] = row1_data[239] ? 16'b0 : row1_data[239:224];
    assign act_row1_data[255:240] = row1_data[255] ? 16'b0 : row1_data[255:240];

    assign act_row2_vld = {16{act_vld}};

    assign act_row2_data[15:0] = row2_data[15] ? 16'b0 : row2_data[15:0];
    assign act_row2_data[31:16] = row2_data[31] ? 16'b0 : row2_data[31:16];
    assign act_row2_data[47:32] = row2_data[47] ? 16'b0 : row2_data[47:32];
    assign act_row2_data[63:48] = row2_data[63] ? 16'b0 : row2_data[63:48];
    assign act_row2_data[79:64] = row2_data[79] ? 16'b0 : row2_data[79:64];
    assign act_row2_data[95:80] = row2_data[95] ? 16'b0 : row2_data[95:80];
    assign act_row2_data[111:96] = row2_data[111] ? 16'b0 : row2_data[111:96];
    assign act_row2_data[127:112] = row2_data[127] ? 16'b0 : row2_data[127:112];
    assign act_row2_data[143:128] = row2_data[143] ? 16'b0 : row2_data[143:128];
    assign act_row2_data[159:144] = row2_data[159] ? 16'b0 : row2_data[159:144];
    assign act_row2_data[175:160] = row2_data[175] ? 16'b0 : row2_data[175:160];
    assign act_row2_data[191:176] = row2_data[191] ? 16'b0 : row2_data[191:176];
    assign act_row2_data[207:192] = row2_data[207] ? 16'b0 : row2_data[207:192];
    assign act_row2_data[223:208] = row2_data[223] ? 16'b0 : row2_data[223:208];
    assign act_row2_data[239:224] = row2_data[239] ? 16'b0 : row2_data[239:224];
    assign act_row2_data[255:240] = row2_data[255] ? 16'b0 : row2_data[255:240];

    assign act_row3_vld = {16{act_vld}};

    assign act_row3_data[15:0] = row3_data[15] ? 16'b0 : row3_data[15:0];
    assign act_row3_data[31:16] = row3_data[31] ? 16'b0 : row3_data[31:16];
    assign act_row3_data[47:32] = row3_data[47] ? 16'b0 : row3_data[47:32];
    assign act_row3_data[63:48] = row3_data[63] ? 16'b0 : row3_data[63:48];
    assign act_row3_data[79:64] = row3_data[79] ? 16'b0 : row3_data[79:64];
    assign act_row3_data[95:80] = row3_data[95] ? 16'b0 : row3_data[95:80];
    assign act_row3_data[111:96] = row3_data[111] ? 16'b0 : row3_data[111:96];
    assign act_row3_data[127:112] = row3_data[127] ? 16'b0 : row3_data[127:112];
    assign act_row3_data[143:128] = row3_data[143] ? 16'b0 : row3_data[143:128];
    assign act_row3_data[159:144] = row3_data[159] ? 16'b0 : row3_data[159:144];
    assign act_row3_data[175:160] = row3_data[175] ? 16'b0 : row3_data[175:160];
    assign act_row3_data[191:176] = row3_data[191] ? 16'b0 : row3_data[191:176];
    assign act_row3_data[207:192] = row3_data[207] ? 16'b0 : row3_data[207:192];
    assign act_row3_data[223:208] = row3_data[223] ? 16'b0 : row3_data[223:208];
    assign act_row3_data[239:224] = row3_data[239] ? 16'b0 : row3_data[239:224];
    assign act_row3_data[255:240] = row3_data[255] ? 16'b0 : row3_data[255:240];

    assign act_row4_vld = {16{act_vld}};

    assign act_row4_data[15:0] = row4_data[15] ? 16'b0 : row4_data[15:0];
    assign act_row4_data[31:16] = row4_data[31] ? 16'b0 : row4_data[31:16];
    assign act_row4_data[47:32] = row4_data[47] ? 16'b0 : row4_data[47:32];
    assign act_row4_data[63:48] = row4_data[63] ? 16'b0 : row4_data[63:48];
    assign act_row4_data[79:64] = row4_data[79] ? 16'b0 : row4_data[79:64];
    assign act_row4_data[95:80] = row4_data[95] ? 16'b0 : row4_data[95:80];
    assign act_row4_data[111:96] = row4_data[111] ? 16'b0 : row4_data[111:96];
    assign act_row4_data[127:112] = row4_data[127] ? 16'b0 : row4_data[127:112];
    assign act_row4_data[143:128] = row4_data[143] ? 16'b0 : row4_data[143:128];
    assign act_row4_data[159:144] = row4_data[159] ? 16'b0 : row4_data[159:144];
    assign act_row4_data[175:160] = row4_data[175] ? 16'b0 : row4_data[175:160];
    assign act_row4_data[191:176] = row4_data[191] ? 16'b0 : row4_data[191:176];
    assign act_row4_data[207:192] = row4_data[207] ? 16'b0 : row4_data[207:192];
    assign act_row4_data[223:208] = row4_data[223] ? 16'b0 : row4_data[223:208];
    assign act_row4_data[239:224] = row4_data[239] ? 16'b0 : row4_data[239:224];
    assign act_row4_data[255:240] = row4_data[255] ? 16'b0 : row4_data[255:240];

    assign act_row5_vld = {16{act_vld}};

    assign act_row5_data[15:0] = row5_data[15] ? 16'b0 : row5_data[15:0];
    assign act_row5_data[31:16] = row5_data[31] ? 16'b0 : row5_data[31:16];
    assign act_row5_data[47:32] = row5_data[47] ? 16'b0 : row5_data[47:32];
    assign act_row5_data[63:48] = row5_data[63] ? 16'b0 : row5_data[63:48];
    assign act_row5_data[79:64] = row5_data[79] ? 16'b0 : row5_data[79:64];
    assign act_row5_data[95:80] = row5_data[95] ? 16'b0 : row5_data[95:80];
    assign act_row5_data[111:96] = row5_data[111] ? 16'b0 : row5_data[111:96];
    assign act_row5_data[127:112] = row5_data[127] ? 16'b0 : row5_data[127:112];
    assign act_row5_data[143:128] = row5_data[143] ? 16'b0 : row5_data[143:128];
    assign act_row5_data[159:144] = row5_data[159] ? 16'b0 : row5_data[159:144];
    assign act_row5_data[175:160] = row5_data[175] ? 16'b0 : row5_data[175:160];
    assign act_row5_data[191:176] = row5_data[191] ? 16'b0 : row5_data[191:176];
    assign act_row5_data[207:192] = row5_data[207] ? 16'b0 : row5_data[207:192];
    assign act_row5_data[223:208] = row5_data[223] ? 16'b0 : row5_data[223:208];
    assign act_row5_data[239:224] = row5_data[239] ? 16'b0 : row5_data[239:224];
    assign act_row5_data[255:240] = row5_data[255] ? 16'b0 : row5_data[255:240];

    assign act_row6_vld = {16{act_vld}};

    assign act_row6_data[15:0] = row6_data[15] ? 16'b0 : row6_data[15:0];
    assign act_row6_data[31:16] = row6_data[31] ? 16'b0 : row6_data[31:16];
    assign act_row6_data[47:32] = row6_data[47] ? 16'b0 : row6_data[47:32];
    assign act_row6_data[63:48] = row6_data[63] ? 16'b0 : row6_data[63:48];
    assign act_row6_data[79:64] = row6_data[79] ? 16'b0 : row6_data[79:64];
    assign act_row6_data[95:80] = row6_data[95] ? 16'b0 : row6_data[95:80];
    assign act_row6_data[111:96] = row6_data[111] ? 16'b0 : row6_data[111:96];
    assign act_row6_data[127:112] = row6_data[127] ? 16'b0 : row6_data[127:112];
    assign act_row6_data[143:128] = row6_data[143] ? 16'b0 : row6_data[143:128];
    assign act_row6_data[159:144] = row6_data[159] ? 16'b0 : row6_data[159:144];
    assign act_row6_data[175:160] = row6_data[175] ? 16'b0 : row6_data[175:160];
    assign act_row6_data[191:176] = row6_data[191] ? 16'b0 : row6_data[191:176];
    assign act_row6_data[207:192] = row6_data[207] ? 16'b0 : row6_data[207:192];
    assign act_row6_data[223:208] = row6_data[223] ? 16'b0 : row6_data[223:208];
    assign act_row6_data[239:224] = row6_data[239] ? 16'b0 : row6_data[239:224];
    assign act_row6_data[255:240] = row6_data[255] ? 16'b0 : row6_data[255:240];

    assign act_row7_vld = {16{act_vld}};

    assign act_row7_data[15:0] = row7_data[15] ? 16'b0 : row7_data[15:0];
    assign act_row7_data[31:16] = row7_data[31] ? 16'b0 : row7_data[31:16];
    assign act_row7_data[47:32] = row7_data[47] ? 16'b0 : row7_data[47:32];
    assign act_row7_data[63:48] = row7_data[63] ? 16'b0 : row7_data[63:48];
    assign act_row7_data[79:64] = row7_data[79] ? 16'b0 : row7_data[79:64];
    assign act_row7_data[95:80] = row7_data[95] ? 16'b0 : row7_data[95:80];
    assign act_row7_data[111:96] = row7_data[111] ? 16'b0 : row7_data[111:96];
    assign act_row7_data[127:112] = row7_data[127] ? 16'b0 : row7_data[127:112];
    assign act_row7_data[143:128] = row7_data[143] ? 16'b0 : row7_data[143:128];
    assign act_row7_data[159:144] = row7_data[159] ? 16'b0 : row7_data[159:144];
    assign act_row7_data[175:160] = row7_data[175] ? 16'b0 : row7_data[175:160];
    assign act_row7_data[191:176] = row7_data[191] ? 16'b0 : row7_data[191:176];
    assign act_row7_data[207:192] = row7_data[207] ? 16'b0 : row7_data[207:192];
    assign act_row7_data[223:208] = row7_data[223] ? 16'b0 : row7_data[223:208];
    assign act_row7_data[239:224] = row7_data[239] ? 16'b0 : row7_data[239:224];
    assign act_row7_data[255:240] = row7_data[255] ? 16'b0 : row7_data[255:240];

    assign act_row8_vld = {16{act_vld}};

    assign act_row8_data[15:0] = row8_data[15] ? 16'b0 : row8_data[15:0];
    assign act_row8_data[31:16] = row8_data[31] ? 16'b0 : row8_data[31:16];
    assign act_row8_data[47:32] = row8_data[47] ? 16'b0 : row8_data[47:32];
    assign act_row8_data[63:48] = row8_data[63] ? 16'b0 : row8_data[63:48];
    assign act_row8_data[79:64] = row8_data[79] ? 16'b0 : row8_data[79:64];
    assign act_row8_data[95:80] = row8_data[95] ? 16'b0 : row8_data[95:80];
    assign act_row8_data[111:96] = row8_data[111] ? 16'b0 : row8_data[111:96];
    assign act_row8_data[127:112] = row8_data[127] ? 16'b0 : row8_data[127:112];
    assign act_row8_data[143:128] = row8_data[143] ? 16'b0 : row8_data[143:128];
    assign act_row8_data[159:144] = row8_data[159] ? 16'b0 : row8_data[159:144];
    assign act_row8_data[175:160] = row8_data[175] ? 16'b0 : row8_data[175:160];
    assign act_row8_data[191:176] = row8_data[191] ? 16'b0 : row8_data[191:176];
    assign act_row8_data[207:192] = row8_data[207] ? 16'b0 : row8_data[207:192];
    assign act_row8_data[223:208] = row8_data[223] ? 16'b0 : row8_data[223:208];
    assign act_row8_data[239:224] = row8_data[239] ? 16'b0 : row8_data[239:224];
    assign act_row8_data[255:240] = row8_data[255] ? 16'b0 : row8_data[255:240];

    assign act_row9_vld = {16{act_vld}};

    assign act_row9_data[15:0] = row9_data[15] ? 16'b0 : row9_data[15:0];
    assign act_row9_data[31:16] = row9_data[31] ? 16'b0 : row9_data[31:16];
    assign act_row9_data[47:32] = row9_data[47] ? 16'b0 : row9_data[47:32];
    assign act_row9_data[63:48] = row9_data[63] ? 16'b0 : row9_data[63:48];
    assign act_row9_data[79:64] = row9_data[79] ? 16'b0 : row9_data[79:64];
    assign act_row9_data[95:80] = row9_data[95] ? 16'b0 : row9_data[95:80];
    assign act_row9_data[111:96] = row9_data[111] ? 16'b0 : row9_data[111:96];
    assign act_row9_data[127:112] = row9_data[127] ? 16'b0 : row9_data[127:112];
    assign act_row9_data[143:128] = row9_data[143] ? 16'b0 : row9_data[143:128];
    assign act_row9_data[159:144] = row9_data[159] ? 16'b0 : row9_data[159:144];
    assign act_row9_data[175:160] = row9_data[175] ? 16'b0 : row9_data[175:160];
    assign act_row9_data[191:176] = row9_data[191] ? 16'b0 : row9_data[191:176];
    assign act_row9_data[207:192] = row9_data[207] ? 16'b0 : row9_data[207:192];
    assign act_row9_data[223:208] = row9_data[223] ? 16'b0 : row9_data[223:208];
    assign act_row9_data[239:224] = row9_data[239] ? 16'b0 : row9_data[239:224];
    assign act_row9_data[255:240] = row9_data[255] ? 16'b0 : row9_data[255:240];

    assign act_row10_vld = {16{act_vld}};

    assign act_row10_data[15:0] = row10_data[15] ? 16'b0 : row10_data[15:0];
    assign act_row10_data[31:16] = row10_data[31] ? 16'b0 : row10_data[31:16];
    assign act_row10_data[47:32] = row10_data[47] ? 16'b0 : row10_data[47:32];
    assign act_row10_data[63:48] = row10_data[63] ? 16'b0 : row10_data[63:48];
    assign act_row10_data[79:64] = row10_data[79] ? 16'b0 : row10_data[79:64];
    assign act_row10_data[95:80] = row10_data[95] ? 16'b0 : row10_data[95:80];
    assign act_row10_data[111:96] = row10_data[111] ? 16'b0 : row10_data[111:96];
    assign act_row10_data[127:112] = row10_data[127] ? 16'b0 : row10_data[127:112];
    assign act_row10_data[143:128] = row10_data[143] ? 16'b0 : row10_data[143:128];
    assign act_row10_data[159:144] = row10_data[159] ? 16'b0 : row10_data[159:144];
    assign act_row10_data[175:160] = row10_data[175] ? 16'b0 : row10_data[175:160];
    assign act_row10_data[191:176] = row10_data[191] ? 16'b0 : row10_data[191:176];
    assign act_row10_data[207:192] = row10_data[207] ? 16'b0 : row10_data[207:192];
    assign act_row10_data[223:208] = row10_data[223] ? 16'b0 : row10_data[223:208];
    assign act_row10_data[239:224] = row10_data[239] ? 16'b0 : row10_data[239:224];
    assign act_row10_data[255:240] = row10_data[255] ? 16'b0 : row10_data[255:240];

    assign act_row11_vld = {16{act_vld}};

    assign act_row11_data[15:0] = row11_data[15] ? 16'b0 : row11_data[15:0];
    assign act_row11_data[31:16] = row11_data[31] ? 16'b0 : row11_data[31:16];
    assign act_row11_data[47:32] = row11_data[47] ? 16'b0 : row11_data[47:32];
    assign act_row11_data[63:48] = row11_data[63] ? 16'b0 : row11_data[63:48];
    assign act_row11_data[79:64] = row11_data[79] ? 16'b0 : row11_data[79:64];
    assign act_row11_data[95:80] = row11_data[95] ? 16'b0 : row11_data[95:80];
    assign act_row11_data[111:96] = row11_data[111] ? 16'b0 : row11_data[111:96];
    assign act_row11_data[127:112] = row11_data[127] ? 16'b0 : row11_data[127:112];
    assign act_row11_data[143:128] = row11_data[143] ? 16'b0 : row11_data[143:128];
    assign act_row11_data[159:144] = row11_data[159] ? 16'b0 : row11_data[159:144];
    assign act_row11_data[175:160] = row11_data[175] ? 16'b0 : row11_data[175:160];
    assign act_row11_data[191:176] = row11_data[191] ? 16'b0 : row11_data[191:176];
    assign act_row11_data[207:192] = row11_data[207] ? 16'b0 : row11_data[207:192];
    assign act_row11_data[223:208] = row11_data[223] ? 16'b0 : row11_data[223:208];
    assign act_row11_data[239:224] = row11_data[239] ? 16'b0 : row11_data[239:224];
    assign act_row11_data[255:240] = row11_data[255] ? 16'b0 : row11_data[255:240];

    assign act_row12_vld = {16{act_vld}};

    assign act_row12_data[15:0] = row12_data[15] ? 16'b0 : row12_data[15:0];
    assign act_row12_data[31:16] = row12_data[31] ? 16'b0 : row12_data[31:16];
    assign act_row12_data[47:32] = row12_data[47] ? 16'b0 : row12_data[47:32];
    assign act_row12_data[63:48] = row12_data[63] ? 16'b0 : row12_data[63:48];
    assign act_row12_data[79:64] = row12_data[79] ? 16'b0 : row12_data[79:64];
    assign act_row12_data[95:80] = row12_data[95] ? 16'b0 : row12_data[95:80];
    assign act_row12_data[111:96] = row12_data[111] ? 16'b0 : row12_data[111:96];
    assign act_row12_data[127:112] = row12_data[127] ? 16'b0 : row12_data[127:112];
    assign act_row12_data[143:128] = row12_data[143] ? 16'b0 : row12_data[143:128];
    assign act_row12_data[159:144] = row12_data[159] ? 16'b0 : row12_data[159:144];
    assign act_row12_data[175:160] = row12_data[175] ? 16'b0 : row12_data[175:160];
    assign act_row12_data[191:176] = row12_data[191] ? 16'b0 : row12_data[191:176];
    assign act_row12_data[207:192] = row12_data[207] ? 16'b0 : row12_data[207:192];
    assign act_row12_data[223:208] = row12_data[223] ? 16'b0 : row12_data[223:208];
    assign act_row12_data[239:224] = row12_data[239] ? 16'b0 : row12_data[239:224];
    assign act_row12_data[255:240] = row12_data[255] ? 16'b0 : row12_data[255:240];

    assign act_row13_vld = {16{act_vld}};

    assign act_row13_data[15:0] = row13_data[15] ? 16'b0 : row13_data[15:0];
    assign act_row13_data[31:16] = row13_data[31] ? 16'b0 : row13_data[31:16];
    assign act_row13_data[47:32] = row13_data[47] ? 16'b0 : row13_data[47:32];
    assign act_row13_data[63:48] = row13_data[63] ? 16'b0 : row13_data[63:48];
    assign act_row13_data[79:64] = row13_data[79] ? 16'b0 : row13_data[79:64];
    assign act_row13_data[95:80] = row13_data[95] ? 16'b0 : row13_data[95:80];
    assign act_row13_data[111:96] = row13_data[111] ? 16'b0 : row13_data[111:96];
    assign act_row13_data[127:112] = row13_data[127] ? 16'b0 : row13_data[127:112];
    assign act_row13_data[143:128] = row13_data[143] ? 16'b0 : row13_data[143:128];
    assign act_row13_data[159:144] = row13_data[159] ? 16'b0 : row13_data[159:144];
    assign act_row13_data[175:160] = row13_data[175] ? 16'b0 : row13_data[175:160];
    assign act_row13_data[191:176] = row13_data[191] ? 16'b0 : row13_data[191:176];
    assign act_row13_data[207:192] = row13_data[207] ? 16'b0 : row13_data[207:192];
    assign act_row13_data[223:208] = row13_data[223] ? 16'b0 : row13_data[223:208];
    assign act_row13_data[239:224] = row13_data[239] ? 16'b0 : row13_data[239:224];
    assign act_row13_data[255:240] = row13_data[255] ? 16'b0 : row13_data[255:240];

    assign act_row14_vld = {16{act_vld}};

    assign act_row14_data[15:0] = row14_data[15] ? 16'b0 : row14_data[15:0];
    assign act_row14_data[31:16] = row14_data[31] ? 16'b0 : row14_data[31:16];
    assign act_row14_data[47:32] = row14_data[47] ? 16'b0 : row14_data[47:32];
    assign act_row14_data[63:48] = row14_data[63] ? 16'b0 : row14_data[63:48];
    assign act_row14_data[79:64] = row14_data[79] ? 16'b0 : row14_data[79:64];
    assign act_row14_data[95:80] = row14_data[95] ? 16'b0 : row14_data[95:80];
    assign act_row14_data[111:96] = row14_data[111] ? 16'b0 : row14_data[111:96];
    assign act_row14_data[127:112] = row14_data[127] ? 16'b0 : row14_data[127:112];
    assign act_row14_data[143:128] = row14_data[143] ? 16'b0 : row14_data[143:128];
    assign act_row14_data[159:144] = row14_data[159] ? 16'b0 : row14_data[159:144];
    assign act_row14_data[175:160] = row14_data[175] ? 16'b0 : row14_data[175:160];
    assign act_row14_data[191:176] = row14_data[191] ? 16'b0 : row14_data[191:176];
    assign act_row14_data[207:192] = row14_data[207] ? 16'b0 : row14_data[207:192];
    assign act_row14_data[223:208] = row14_data[223] ? 16'b0 : row14_data[223:208];
    assign act_row14_data[239:224] = row14_data[239] ? 16'b0 : row14_data[239:224];
    assign act_row14_data[255:240] = row14_data[255] ? 16'b0 : row14_data[255:240];

    assign act_row15_vld = {16{act_vld}};

    assign act_row15_data[15:0] = row15_data[15] ? 16'b0 : row15_data[15:0];
    assign act_row15_data[31:16] = row15_data[31] ? 16'b0 : row15_data[31:16];
    assign act_row15_data[47:32] = row15_data[47] ? 16'b0 : row15_data[47:32];
    assign act_row15_data[63:48] = row15_data[63] ? 16'b0 : row15_data[63:48];
    assign act_row15_data[79:64] = row15_data[79] ? 16'b0 : row15_data[79:64];
    assign act_row15_data[95:80] = row15_data[95] ? 16'b0 : row15_data[95:80];
    assign act_row15_data[111:96] = row15_data[111] ? 16'b0 : row15_data[111:96];
    assign act_row15_data[127:112] = row15_data[127] ? 16'b0 : row15_data[127:112];
    assign act_row15_data[143:128] = row15_data[143] ? 16'b0 : row15_data[143:128];
    assign act_row15_data[159:144] = row15_data[159] ? 16'b0 : row15_data[159:144];
    assign act_row15_data[175:160] = row15_data[175] ? 16'b0 : row15_data[175:160];
    assign act_row15_data[191:176] = row15_data[191] ? 16'b0 : row15_data[191:176];
    assign act_row15_data[207:192] = row15_data[207] ? 16'b0 : row15_data[207:192];
    assign act_row15_data[223:208] = row15_data[223] ? 16'b0 : row15_data[223:208];
    assign act_row15_data[239:224] = row15_data[239] ? 16'b0 : row15_data[239:224];
    assign act_row15_data[255:240] = row15_data[255] ? 16'b0 : row15_data[255:240];


endmodule 