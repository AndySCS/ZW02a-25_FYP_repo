import uvm_pkg::*;