python3 ../regression/regression.py --list ../regression/regression_list.json
