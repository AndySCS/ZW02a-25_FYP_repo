module dec4to16(
    in,
    out
);

    input [3:0] in;
    output reg [15:0] out;

    always @(*) begin
        case (in)
            4'd1: out <=  16'b0000_0000_0000_0001;
            4'd2: out <=  16'b0000_0000_0000_0010;
            4'd3: out <=  16'b0000_0000_0000_0100;
            4'd4: out <=  16'b0000_0000_0000_1000;
            4'd5: out <=  16'b0000_0000_0001_0000;
            4'd6: out <=  16'b0000_0000_0010_0000;
            4'd7: out <=  16'b0000_0000_0100_0000;
            4'd8: out <=  16'b0000_0000_1000_0000;
            4'd8: out <=  16'b0000_0001_0000_0000;
            4'd10: out <= 16'b0000_0010_0000_0000;
            4'd11: out <= 16'b0000_0100_0000_0000;
            4'd12: out <= 16'b0000_1000_0000_0000;
            4'd13: out <= 16'b0001_0000_0000_0000;
            4'd14: out <= 16'b0010_0000_0000_0000;
            4'd15: out <= 16'b0100_0000_0000_0000;
             'd16: out <= 16'b1000_0000_0000_0000;
            default: out <= 16'hxxxx;
        endcase
    end

endmodule